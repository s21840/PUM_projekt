��}�      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �min_impurity_split�N�class_weight�N�	ccp_alpha�G        �_sklearn_version��0.24.2�ub�n_estimators�K�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK�verbose�K �
warm_start��hN�max_samples�NhhhKhKhKhG        h�auto�hNhG        hNhG        �n_features_in_�K�n_features_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h-�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhKhKhKhG        hh%hNhJc��8hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��h6�f8�����R�(Kh:NNNJ����J����K t�b�C              �?�t�bh>h*�scalar���h9C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hK�
node_count�K��nodes�h,h/K ��h1��R�(KK���h6�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hkh9K ��hlh9K��hmh9K��hnhJK��hohJK ��hph9K(��hqhJK0��uK8KKt�b�BX"         6                 � >濂sF����?�           @�@                        0���?l��(��?6           ��@                        �0	�?�:��?k           ��@                         0�M�?���.I��?=           ��@������������������������       �                   @�@       	                 нA�h�WH��?              K@                        0_�? ���J��?            �C@������������������������       �                     C@������������������������       �                     �?
                        PY�ῲ�����?	             .@������������������������       �                      @                         ���?8�Z$���?             *@������������������������       �                     @                         ����?����X�?             @������������������������       �                      @������������������������       �                     @                        `G��? � {�o?.           0�@������������������������       �        *            �@                        �;��?r�q��?             @������������������������       �                     �?������������������������       �                     @       5                 �Z��?|��?���?�            @t@       2                 �0	�?\x�R:��?�            Ps@       +                 P��Ŀ���7ۨ�?�            �k@                         �J�ۿ��=A��?1             S@������������������������       �                     8@       *                 p4�?���c���?"             J@                        P@�?fP*L��?             F@                        ��1�?���|���?             &@������������������������       �                     @������������������������       �                     @        !                 @6`�?�C��2(�?            �@@������������������������       �                     1@"       %                 0�8ƿ     ��?
             0@#       $                  @���?���Q��?             @������������������������       �                     @������������������������       �                      @&       '                 ��uſ�C��2(�?             &@������������������������       �                     @(       )                 �Xcſz�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @,       1                 p4�?�Q���?\            `b@-       .                 ��Z�t�0i��?W            `a@������������������������       �        &             L@/       0                  �3�?�L"p�?1            �T@������������������������       �                    �G@������������������������       �                     B@������������������������       �                      @3       4                  H=�?8�$�>�?3            �U@������������������������       �                      L@������������������������       �                     >@������������������������       �                     .@7       ~                 p4�?& ����?]           X�@8       ]                 �0	�?~�ӻH��?�           �@9       \                 �Ƴ�?�ήxF�?V
           H�@:       =                 ��Z󿾺i�?�	           ��@;       <                  �ˑ?~|z����?�            0w@������������������������       �        s            �e@������������������������       �                    �h@>       [                  �� �?�@��*��?�           ث@?       T                  ��?NW����?�           �@@       O                 �P�?ޝ8t|}�?           0�@A       J                  ��k�?��f�?�           ޢ@B       C                 �8�ƿ,���-v�?�           ��@������������������������       �                     "@D       G                  0�IۿJ
{�}�?�           ��@E       F                 �pm¿~���L0�?_            `b@������������������������       ��le����?A            �Z@������������������������       ��Q����?             D@H       I                 ����?&��F��?�           t�@������������������������       �        ~           �@������������������������       �                   \�@K       L                 �tƿHP�s��?             9@������������������������       �                     �?M       N                 ���ο �q�q�?             8@������������������������       �                     �?������������������������       �                     7@P       Q                 ����?���?            �D@������������������������       �                     .@R       S                 p��ȿ�n_Y�K�?             :@������������������������       �                     0@������������������������       �                     $@U       X                 ��?�|�a�B�?�             k@V       W                 ��`�?�kwY���?�            @j@������������������������       �        G             _@������������������������       �        9            �U@Y       Z                 	J�?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        @           ؋@������������������������       �        �             m@^       q                  ���?z��=��?<           P�@_       b                  @ҙ��h��ݥ��?$           ��@`       a                 �
��?ܥ8Pj{�?Q            �@������������������������       �        n           p�@������������������������       �        �           Ї@c       f                 �mĿF��ӭ��?�            �v@d       e                 @[M�?&��QK?�?d            `d@������������������������       �        +            @Q@������������������������       �        9            �W@g       j                  �ÿ�1׹k��?o            �h@h       i                 ����?"pc�
�?             F@������������������������       �                     B@������������������������       �                      @k       n                  �4<�?N�[7���?W             c@l       m                 @�+���û��|�?4             W@������������������������       �                     L@������������������������       �                     B@o       p                  5�z?�u���?#            �N@������������������������       �                     8@������������������������       �                    �B@r       y                  ��^��4?,R��?             B@s       x                  �#�ӿףp=
�?             >@t       u                 ��Z�@�0�!��?             1@������������������������       �                      @v       w                 @�V���q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     *@z       }                 P��@�q�q�?             @{       |                  �w�?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?       �                  �s\�?p��D׀�?�            �s@�       �                 @^�? %��$��?�            r@�       �                 �:��?�s�}?�            �q@������������������������       �        �             q@�       �                 p| �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                  0��ڿ      �?              @������������������������       �                     @������������������������       �                     @�       �                 ��qƿ|��?���?             ;@�       �                  1���z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                 0]�ſ�eP*L��?             6@�       �                 Pt/ƿ؇���X�?             @������������������������       �                     @�       �                 X�&�?      �?             @������������������������       �                     @������������������������       �                     �?�       �                  �*	�?���Q��?             .@�       �                 p�nƿ      �?              @������������������������       �                     �?������������������������       �                     @�       �                  `��?����X�?             @������������������������       �                     @�       �                 �0	�?      �?             @�       �                  �=o?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�t�b�values�h,h/K ��h1��R�(KK�KK��hJ�B�	       ��@     �@     �@     �e@     x�@      @     Ȍ@      @     @�@             �H@      @      C@      �?      C@                      �?      &@      @               @      &@       @      @              @       @               @      @             (�@      �?      �@              @      �?              �?      @             �c@      e@     �c@      c@      Y@     �^@     �F@      ?@              8@     �F@      @     �B@      @      @      @      @                      @      >@      @      1@              *@      @      @       @      @                       @      $@      �?      @              @      �?              �?      @               @             �K@      W@     �G@      W@              L@     �G@      B@     �G@                      B@       @              L@      >@      L@                      >@              .@     &�@     ��@     Ҡ@     f�@     t�@     ֥@     t�@     �@     �e@     �h@     �e@                     �h@     ��@     |�@     ��@     �@     Đ@     ��@     H�@     t�@     @�@     �@              "@     @�@     ��@     �F@     �Y@      :@     @T@      3@      5@     �@     \�@     �@                     \�@       @      7@      �?              �?      7@      �?                      7@      ?@      $@      .@              0@      $@      0@                      $@     @_@      W@      _@     �U@      _@                     �U@      �?      @              @      �?                     ؋@              m@     `�@     @�@     8�@     H�@     p�@     Ї@     p�@                     Ї@      g@     �e@     @Q@     �W@     @Q@                     �W@      ]@     @T@      B@       @      B@                       @      T@     @R@      L@      B@      L@                      B@      8@     �B@      8@                     �B@      @      ?@      @      ;@      @      ,@               @      @      @      @                      @              *@       @      @      �?      @      �?                      @      �?             �r@      2@     �q@      @     �q@      �?      q@              @      �?      @                      �?      @      @              @      @              *@      ,@      �?      @      �?                      @      (@      $@      @      �?      @              @      �?      @                      �?      @      "@      �?      @      �?                      @      @       @      @               @       @      �?       @      �?                       @      �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh%hNhJ�H hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaKuhbh,h/K ��h1��R�(KKu��hi�B�         P                  �h
�?N|��8��?�           @�@       I                 p4�?�F���D�?�           }�@       "                 �ʑ�?h�Q�?�           ��@                         Ķ�?��˒5J�?�           ̫@������������������������       �        ;           ��@                        @���?4�dS���?�            pp@                          �VͿ��}���?4            @S@       	                 ���⿀X�<ݺ?%             K@������������������������       �                     8@
                        ��R�ףp=
�?             >@������������������������       �                     �?                        �0	�? 	��p�?             =@������������������������       �                     ;@������������������������       �                      @                        � >�8����?             7@������������������������       �                     @                        @��翈IєX�?             1@������������������������       �                     �?������������������������       �                     0@                        � >� rpa�?v            @g@������������������������       �                     @                        ��6#@�&���?s            �f@                        �0	�?��Bs�?n            �e@������������������������       �        e            �c@                        �}�?     ��?	             0@������������������������       �                     @                         ����z�G��?             $@������������������������       �                     @                        �1��?���Q��?             @������������������������       �                     @������������������������       �                      @        !                  �[)@      �?              @������������������������       �                      @������������������������       �                     @#       &                 ��ֱ?��;V7��?�           ��@$       %                 � >濲�����?             .@������������������������       �                     @������������������������       �                     &@'       H                 � >��A�.�?�           ~�@(       ;                 ��Z󿠸)���?�             m@)       ,                 @��ƿh�V���?>             V@*       +                 �n��?�q�q�?             @������������������������       �                     �?������������������������       �                      @-       4                   Ãܿ�m(�X�?<            @U@.       /                 ����?@�0�!��?	             1@������������������������       �                      @0       3                  �ܿ��S�ۿ?             .@1       2                 � ��?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@5       8                  -S���IєX�?3             Q@6       7                 �0	�?h�����?*             L@������������������������       �        (             K@������������������������       �                      @9       :                 �)���r�q��?	             (@������������������������       �                      @������������������������       �                     $@<       ?                  `�ֿ֦:O���?X             b@=       >                 t�L�?�i�y�?&            �O@������������������������       �        %            �N@������������������������       �                      @@       C                 �0	�?���� �?2            �T@A       B                 0ʓ�?&y�X���?$             M@������������������������       �                    �G@������������������������       �                     &@D       E                 p5��?r�q��?             8@������������������������       �                     @F       G                  @�E˿��Q��?             4@������������������������       �                     @������������������������       �                     *@������������������������       �        1           ��@J       K                 � >��]J�>��?'           �|@������������������������       �        l             e@L       M                 0�V�?�"��	�?�            r@������������������������       �        �            �q@N       O                 (���?      �?              @������������������������       �                     @������������������������       �                     @Q       `                 �0	�?<�:��_�?           �@R       [                 p4�?�ӖF2��?�           ��@S       Z                 � >濸�GeϹ?�           $�@T       Y                 `w����7i���?>            �Y@U       X                  �J@     ��?%             P@V       W                 Ы��?X��Oԣ�?$             O@������������������������       �                     �K@������������������������       �                     @������������������������       �                      @������������������������       �                     C@������������������������       �        Q           �@\       _                  �>@      �?             @@]       ^                 `E��?8^s]e�?             =@������������������������       �                     4@������������������������       �                     "@������������������������       �                     @a       t                 p4�?�J��?b            @c@b       o                 � >�$ m���?[            @b@c       h                   X��?�w��#��?!             I@d       e                  `�~�?�	j*D�?             *@������������������������       �                     �?f       g                  {]�      �?             (@������������������������       �                     "@������������������������       �                     @i       n                 �ٿ���@��?            �B@j       k                  F��?�����H�?             "@������������������������       �                     @l       m                 �_��z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     <@p       s                ���¢?      �?:             X@q       r                 �`��?�}�+r��?             C@������������������������       �                     B@������������������������       �                      @������������������������       �        !             M@������������������������       �                      @�t�bh~h,h/K ��h1��R�(KKuKK��hJ�BP       ��@     �@     ~�@     |�@     �@     v�@     �@     `n@     ��@              4@     `n@      $@     �P@      @     �I@              8@      @      ;@      �?               @      ;@              ;@       @              @      0@      @              �?      0@      �?                      0@      $@      f@      @              @      f@      @     @e@             �c@      @      *@              @      @      @              @      @       @      @                       @       @      @       @                      @     �`@     ��@      @      &@      @                      &@     @`@     z�@     @`@     �Y@      "@     �S@       @      �?              �?       @              @     �S@      @      ,@       @              �?      ,@      �?      @      �?                      @              $@      @      P@       @      K@              K@       @               @      $@       @                      $@     @^@      8@     �N@       @     �N@                       @      N@      6@     �G@      &@     �G@                      &@      *@      &@              @      *@      @              @      *@                     ��@     `|@      @      e@             �q@      @     �q@              @      @              @      @              a@     �@     �R@     ��@     �K@     ��@     �K@     �G@     �K@      "@     �K@      @     �K@                      @               @              C@             �@      4@      (@      4@      "@      4@                      "@              @     �N@     @W@     �J@     @W@      1@     �@@      "@      @              �?      "@      @      "@                      @       @      =@       @      �?      @              @      �?              �?      @                      <@      B@      N@      B@       @      B@                       @              M@       @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh%hNhJ�O�^hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hK
haKohbh,h/K ��h1��R�(KKo��hi�BH         (                 � >�&���L��?�           @�@                        08�?L��� �?/           |�@                        ��Z� �e���q?c           l�@������������������������       �        i            �d@                        P��翀�Ʈ�Ot?�           ܒ@       	                 �0	�? 7���B�?             K@                        �v��?�(\����?             D@������������������������       �                    �C@������������������������       �                     �?
                         `���?@4և���?             ,@������������������������       �                     *@������������������������       �                     �?                        ����? :|�&e\?�           �@������������������������       �        �           �@                         İ��?؇���X�?             @������������������������       �                     @������������������������       �                     �?       !                 ��Z�(Q��h�?�            @t@                         P��ۿ�*v��?A            @X@                        ����?�nkK�?=             W@                        �0	�?      �?             (@������������������������       �                     "@������������������������       �                     @                         `��ܿ@�z�G�?5             T@                        ps��?      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �        /             R@                        0j4�?���Q��?             @������������������������       �                      @                         ��ſ�q�q�?             @������������������������       �                     �?������������������������       �                      @"       '                  h�w�?�������?�            `l@#       &                 p4�?�����?]            �b@$       %                 pHm�?�5̾�?P            �_@������������������������       �        G            @\@������������������������       �        	             ,@������������������������       �                     5@������������������������       �        .            �S@)       R                 0�?r�<���?�           ��@*       1                  -r�? J��2 �?�           ��@+       ,                  @6��?�7���?           �@������������������������       �        �            �@-       0                 p4�?P��t�x�?$           �@.       /                 �0	�?ptk$�P�?           H�@������������������������       �                   �@������������������������       �                     C@������������������������       �                     8@2       C                 ��P�?��{��w�?�           *�@3       4                 p4�?�������?^           �@������������������������       �        F           ��@5       B                 �0	�?�\��N��?             C@6       =                 �)Ŀ��
P��?            �A@7       <                  ��Ŀ���!pc�?             6@8       ;                 p���?��
ц��?	             *@9       :                  ��Q�?���|���?             &@������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     "@>       ?                 p����8�Z$���?             *@������������������������       �                     @@       A                  �O��?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @D       G                 ��Z���(-�?`            @b@E       F                 p4�?z�G�z�?             $@������������������������       �                      @������������������������       �                      @H       O                 `7a�?г�wY;�?Y             a@I       N                 �0	�?��a�n`�?             ?@J       M                  ~�?R���Q�?             4@K       L                 `x�?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �        	             ,@������������������������       �                     &@P       Q                 p4�?@��!�Q�?E            @Z@������������������������       �        D             Z@������������������������       �                     �?S       T                 ��Z�X;��?�            �p@������������������������       �                     A@U       h                 `�>@�)�9N�?�             m@V       c                 p4�? ��>χ�?�             k@W       \                 `6�翠ջ����?�             j@X       [                 ����?      �?              @Y       Z                 �0	�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @]       b                 "\�?@��d�`�?�             i@^       a                 p��ٿףp=
�?             $@_       `                 �0	�?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        |            �g@d       g                 �� @X�<ݚ�?             "@e       f                  ��-ڿ�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @i       n                  �`�?     ��?             0@j       m                  ���ֿ@4և���?             ,@k       l                 �$@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�t�bh~h,h/K ��h1��R�(KKoKK��hJ�B�       ��@     ��@     ��@     `g@     `�@      @     �d@             В@      @      J@       @     �C@      �?     �C@                      �?      *@      �?      *@                      �?      �@      �?     �@              @      �?      @                      �?     �a@      g@      @     �V@      @      V@      @      "@              "@      @              �?     �S@      �?      @      �?                      @              R@       @      @               @       @      �?              �?       @             �`@     @W@     �`@      ,@     @\@      ,@     @\@                      ,@      5@                     �S@     £@     ��@     ��@     |�@     |�@     �@      �@              O@     �@      C@     �@             �@      C@              8@              :@     ��@      4@     ޣ@             ��@      4@      2@      1@      2@      @      0@      @      @      @      @      @                      @       @                      "@      &@       @      @              @       @      @                       @      @              @     �a@       @       @               @       @              @     �`@      @      <@      @      1@      @      @              @      @                      ,@              &@      �?      Z@              Z@      �?              "@      p@              A@      "@      l@      @     `j@       @     �i@      �?      @      �?       @               @      �?                      @      �?     �h@      �?      "@      �?      @              @      �?                      @             �g@      @      @      @       @               @      @                      @      @      *@      �?      *@      �?      @              @      �?                       @       @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh%hNhJ���ThG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B�         t                 p4�?кFˁ��?�           @�@       5                  q�?�iF@��?e           B�@                        � >��&9���?           ��@                        ��l�? ���v�?           x�@������������������������       �                   ,�@                        ��'޿�\��N��?             3@                        �0	�?      �?	             (@       	                 �T��?�z�G��?             $@������������������������       �                     @
                        `���և���X�?             @������������������������       �                      @                         p�Y�?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @       &                  ���?�6ݔ�1�?�           �@                        �0	�?������?�           @�@                        p��Կ�:pΈ��?�            �@                         ��@ܿħ�/|��?W           �@������������������������       �        &             K@                        ��c�?0��l��?1           8�@������������������������       �        �           |�@������������������������       �        q            �e@                        H���?tk~X��?�            �o@������������������������       �        �            `i@������������������������       �                    �H@       %                 ��Z��û��?�            �@                         �8�濬ܸb���?A             W@                        �  @�z�G��?             $@������������������������       �                     @������������������������       �                     @!       "                 @׎���p\�?<            �T@������������������������       �                     :@#       $                 `���? �Cc}�?*             L@������������������������       �        &             I@������������������������       �                     @������������������������       �        �            �@'       2                  pe��? ��IO�?           ��@(       +                 ����Tc�?x           ��@)       *                 �0	�?hA� �?            �~@������������������������       �                   P}@������������������������       �                     5@,       -                 0'׷?���б�?X            �`@������������������������       �        5            @T@.       /                 �0	�?@3����?#             K@������������������������       �                    �G@0       1                  ���?؇���X�?             @������������������������       �                     �?������������������������       �                     @3       4                 �0	�?�=_���?�            �k@������������������������       �        �            �i@������������������������       �        
             0@6       a                 �.�?�aL�4(�?d           h�@7       `                 � >濰��	���?>           ��@8       C                 ��Z�h �`�?�            `m@9       B                 v��? wVX(6�?-            @T@:       A                 0=*�?L紂P�?            �I@;       <                 �0	�?�8��8��?             H@������������������������       �                     D@=       >                 ���?      �?              @������������������������       �                     @?       @                   ��ۿz�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     >@D       Y                 � ��?8�A�0��?d            @c@E       T                 `-�?Ph�e���?U            �`@F       O                 ��m�?0�n&��?L            �]@G       J                 �0	�?���dQ'�?I            �\@H       I                  �5��?ޚ)�?0             R@������������������������       �                     �G@������������������������       �                     9@K       N                 �v��X�Cc�?             E@L       M                  �N��?�q�q�?             B@������������������������       �                     5@������������������������       �        
             .@������������������������       �                     @P       Q                 ����?z�G�z�?             @������������������������       �                     @R       S                  �K�?      �?              @������������������������       �                     �?������������������������       �                     �?U       V                 �m��?@4և���?	             ,@������������������������       �                     $@W       X                 �2�ƿ      �?             @������������������������       �                     @������������������������       �                     �?Z       [                  ��d��؇���X�?             5@������������������������       �        	             &@\       _                  lW��?�z�G��?             $@]       ^                 �=��?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        �           \�@b       s                 � >激�/�3�?&           ��@c       h                 ��Z�ޚ)�?0             R@d       e                 p�%�?�#-���?            �A@������������������������       �                     7@f       g                 ���ſ      �?             (@������������������������       �                     @������������������������       �                     "@i       l                 ���?�Gi����?            �B@j       k                  � ޱ?b�2�tk�?             2@������������������������       �                     @������������������������       �                     &@m       r                  t���?���y4F�?             3@n       o                 ��@      �?             0@������������������������       �                     &@p       q                 ���	@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        �           P�@u       �                 �0	�?h�|�6�?D           �@v       {                 ��Z�pS0����?�            �w@w       x                 %��?0�)AU��?             �L@������������������������       �                    �J@y       z                  0$8ܿ      �?             @������������������������       �                     @������������������������       �                     �?|       �                  0��?p4�w�?�            �s@}       ~                 @^�?�i��Lg�?�            pr@������������������������       �        �            `q@       �                 4�e�?ҳ�wY;�?	             1@������������������������       �                     &@������������������������       �                     @�       �                 � >��q�q�?             8@������������������������       �                     �?�       �                  Ђ}�?�û��|�?             7@������������������������       �                     $@�       �                 �yſ�	j*D�?	             *@�       �                  �)@؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                 0E���      �?             @������������������������       �                     @������������������������       �                     @������������������������       �        Z            �`@�t�bh~h,h/K ��h1��R�(KK�KK��hJ�B�       ��@     Ԯ@     ګ@     ��@     �@     p�@     T�@      "@     ,�@              $@      "@      @      "@      @      @              @      @      @               @      @       @      @                       @               @      @             ��@     L�@     n�@      m@     ��@      l@     T�@     �e@      K@             |�@     �e@     |�@                     �e@     `i@     �H@     `i@                     �H@     ��@      "@     �T@      "@      @      @      @                      @      S@      @      :@              I@      @      I@                      @      �@              C@     P�@      6@     ؂@      5@     P}@             P}@      5@              �?     �`@             @T@      �?     �J@             �G@      �?      @      �?                      @      0@     �i@             �i@      0@             �^@     r�@     �X@     ��@     �X@      a@      @     �R@      @      F@      @      F@              D@      @      @      @              �?      @      �?                      @      @                      >@     �V@     �O@      V@     �F@     �R@      F@     �R@      D@     �G@      9@     �G@                      9@      ;@      .@      5@      .@      5@                      .@      @              �?      @              @      �?      �?      �?                      �?      *@      �?      $@              @      �?      @                      �?      @      2@              &@      @      @      @      �?      @                      �?              @             \�@      9@     Ȋ@      9@     �G@      @      @@              7@      @      "@      @                      "@      6@      .@      @      &@      @                      &@      .@      @      .@      �?      &@              @      �?              �?      @                      @             P�@     �~@      5@     0v@      5@      L@      �?     �J@              @      �?      @                      �?     �r@      4@     r@      @     `q@              &@      @      &@                      @      $@      ,@      �?              "@      ,@              $@      "@      @      @      �?      @                      �?      @      @              @      @             �`@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh%hNhJ��4hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B�)         �                 
�?8�Վ���?�           @�@                         q�?��\8���?�           ��@                         `��?V�<��o�?�           .�@������������������������       �        )	           �@                        � >��	Ds���?[           X�@������������������������       �        )            �P@                        �0	�?$y�{J��?2           H�@                        ���?���%�?            �@	                        p���� 0?�֎�?�           x�@
                        p4�?@MgzY�?�           p�@������������������������       �        �           (�@������������������������       �                     "@                        �M�ſ�FVQ&�?            �@@                        p4�?      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     9@                        p4�?�����H�?3            @T@������������������������       �        /             R@������������������������       �                     "@������������������������       �                    �D@       )                  @�bۿH�����?G           �@                        � >濐}����?C           �}@                        �0	�?p�eU}�?@            �Y@                         �+�ۿ��F�D�?=            �X@                        p4�?@uvI��?<            �X@������������������������       �        ;            @X@������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       (                 P?��?�m�V_Ʌ?           `w@        %                 0�О���pBI�?3            @R@!       "                  �roۿ@	tbA@�?0            @Q@������������������������       �        -            �P@#       $                 p4�?�q�q�?             @������������������������       �                      @������������������������       �                     �?&       '                  0��ۿ      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        �            �r@*       k                 �0	�?�N^��M�?           J�@+       `                 p4�?$�q-�?�           ��@,       I                 `��?@u���?�           l�@-       0                 @b�ƿ�/a��I�?�           8�@.       /                 � >濶�<b���?             7@������������������������       �                     @������������������������       �                     2@1       H                 � >�p�R]Q�?�           ܒ@2       ;                 pp�?p�|����?A            @\@3       6                 ��Ŀ�GN��?4             V@4       5                  iN �?$�q-�?            �C@������������������������       �                     B@������������������������       �                     @7       :                 �|�n�ڡR����?             �H@8       9                 �ʜ��\X��t�?             G@������������������������       ��&!��?            �E@������������������������       �                     @������������������������       �                     @<       A                 p�|Ŀ� �	��?             9@=       >                 @��?      �?              @������������������������       �                     @?       @                 p�Mƿ      �?             @������������������������       �                     @������������������������       �                     �?B       E                 P?��������?	             1@C       D                 `Ѷ�?$�q-�?             *@������������������������       �                      @������������������������       �z�G�z�?             @F       G                 �&��?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        �           �@J       O                 Y��?�v�ɱ?�            �t@K       N                 � >激��б�?V            �`@L       M                  ��۾?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        R             `@P       U                 |zſ�X�<ݺ?            �h@Q       T                 � >��"w����?1             S@R       S                   ��?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        /            @R@V       W                  h��?85�}C�?N            �^@������������������������       �                     �?X       _                 `;V@\����?M            @^@Y       \                 ��@l��\��?D            �Y@Z       [                 `�j @��<D�m�?A            �X@������������������������       �X�EQ]N�?            �E@������������������������       � �Jj�G�?#            �K@]       ^                  �~@      �?             @������������������������       �                      @������������������������       �      �?              @������������������������       �        	             3@a       j                 �r�?      �?             B@b       i                 �)ĿH�V�e��?             A@c       d                  �>ƿ      �?             ,@������������������������       �                     @e       h                 0��ſ�<ݚ�?             "@f       g                 �3��?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     4@������������������������       �                      @l       u                 ���Ŀ`xA�X�?$           0�@m       t                 � >� ��Q�?�            @x@n       s                 ��:@�X����?             6@o       r                 p4�?      �?             4@p       q                  ����?�E��ӭ�?             2@������������������������       �        	             *@������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �        �            �v@v       �                 @��?���K ]�?7            ~@w       �                 p4�?\TE����?�            `u@x       y                 P��Ŀ�t�5U��?�            �t@������������������������       �                     @z       �                  І�ٿ���Q���?�            �t@{       �                  p��ٿ�S����?"            �L@|                        ��h�?�����H�?              K@}       ~                 � >�      �?             H@������������������������       �                     @������������������������       �                    �F@�       �                 ���?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                 @<��?�I��쪵?�            �p@�       �                 � >�Hb�mS�?�            �p@�       �                 p��?j���� �?             1@������������������������       ����!pc�?             &@������������������������       ��q�q�?             @������������������������       �        �            �o@������������������������       �                      @������������������������       �                     $@�       �                 p4�?P���Q�?X            �a@�       �                  r�@�ㄡ^�?V             a@�       �                  ��6ۿP�c0"�?G            @Z@�       �                 ����?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �        C             Y@�       �                 � >�      �?             @@������������������������       �                      @������������������������       �                     >@������������������������       �                     @�       �                 � >�H%u��?            y@�       �                  P;�ۿNp�����?#            �I@������������������������       �                      @�       �                 p4�?�&!��?            �E@�       �                 �0	�?��%��?            �B@�       �                  ��e�?     ��?             0@�       �                 B�2�?8�Z$���?
             *@������������������������       �                     &@������������������������       �                      @������������������������       �                     @�       �                 �ǳ?և���X�?             5@�       �                   ���?�	j*D�?	             *@������������������������       �                     "@������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                 �0	�?81��=�?�            �u@�       �                 p4�?hڛ�ʚ�?�            �r@�       �                 ��Z󿀃pBI�?�            @r@������������������������       �                    �@@�       �                  ຂۿ`�r��?�            0p@�       �                  �Q�ۿ�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                 ����?     <�?�             p@�       �                 P���?��Q��?             4@�       �                  �XI׿@4և���?             ,@������������������������       �                     �?������������������������       �                     *@������������������������       �                     @������������������������       �        �            �m@�       �                  PN�ؿ�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                 пE߿������?             �I@�       �                 ��Z�      �?             8@������������������������       �                     "@�       �                  �V��?z�G�z�?	             .@������������������������       �                     (@������������������������       �                     @������������������������       �                     ;@�t�bh~h,h/K ��h1��R�(KK�KK��hJ�B�       ܯ@     ��@     |�@     �@     �@     `�@     �@             �_@     `�@     �P@             �N@     `�@      4@     `�@      &@      �@      "@     (�@             (�@      "@               @      ?@       @      @              @       @                      9@      "@      R@              R@      "@             �D@             �g@     ��@       @     P}@      @     @X@       @     @X@      �?     @X@             @X@      �?              �?              @               @     @w@       @     �Q@      �?      Q@             �P@      �?       @               @      �?              �?      @      �?                      @             �r@     �f@     �@     �^@     �@      X@     �@      U@     �@      @      2@      @                      2@     �S@     ��@     �S@      A@     @P@      7@      B@      @      B@                      @      =@      4@      :@      4@      :@      1@              @      @              ,@      &@      �?      @              @      �?      @              @      �?              *@      @      (@      �?       @              @      �?      �?      @              @      �?                     �@      (@     t@      �?     �`@      �?      @      �?                      @              `@      &@     `g@      �?     �R@      �?       @      �?                       @             @R@      $@      \@      �?              "@      \@      "@     @W@      @      W@      @      C@      �?      K@      @      �?       @              �?      �?              3@      ;@      "@      ;@      @      @      @      @               @      @       @      @       @                      @              @      4@                       @     �L@     h�@      .@     Pw@      .@      @      .@      @      *@      @      *@                      @       @                       @             �v@      E@     �{@     �A@     0s@      9@     0s@      @              5@     0s@      "@      H@      @      H@      @     �F@      @                     �F@      @      @      @                      @      @              (@     0p@      $@     0p@      $@      @       @      @       @      @             �o@       @              $@              @     �`@      @     �`@       @     �Y@       @      @       @                      @              Y@       @      >@       @                      >@      @              H@      v@      :@      9@               @      :@      1@      4@      1@      &@      @      &@       @      &@                       @              @      "@      (@      "@      @      "@                      @               @      @              6@     pt@      $@      r@       @     �q@             �@@       @     `o@      �?       @               @      �?              @      o@      @      *@      �?      *@      �?                      *@      @                     �m@       @      @              @       @              (@     �C@      (@      (@              "@      (@      @      (@                      @              ;@�t�bubhhubehhub.