���      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �min_impurity_split�N�class_weight�N�	ccp_alpha�G        �n_features_in_�K�n_features_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�h�scalar���h'C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h'�C       �t�bK��R�}�(h	K�
node_count�K-�nodes�hhK ��h��R�(KK-��h$�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hJh'K ��hKh'K��hLh'K��hMh$�f8�����R�(Kh(NNNJ����J����K t�bK��hNhXK ��hOh'K(��hPhXK0��uK8KKt�b�B�	                          ���@�������?@           @�@                         �i�X@�R��Z�?           �@                        p��H@H��Q6�?^           ��@������������������������       �        O           ��@                           �?	��j�?           �p@������������������������       �                     3@       
                    �?U^C�/��?�            �o@       	                    �?rj�k���?�            �l@������������������������       �        �            �l@������������������������       �                     @                           �?���'���?             5@������������������������       �                     (@������������������������       �        	             "@                           �?5C��Y+�?�           ؍@                        �B�D@|<�;
��?N            �S@������������������������       �        D             Q@������������������������       �        
             $@                           �?�g�����?m           h�@                           �?�r����?B           �@������������������������       �        8           ��@������������������������       �        
             $@                        �aEF@���&��?+            �E@������������������������       �        '            �C@������������������������       �                     @       &                    �?�)Hg���?'           N�@       !                  ��o�?t��#���?X           �u@                           �?i������?t             ]@                           �?'É�,��?o            �[@������������������������       �        m            @[@������������������������       �                      @                         ��B@�Z���?             @������������������������       �                     @������������������������       �                     �?"       %                  ��W@BhBu{E�?�            �l@#       $                 ��GF@_�<��?�            �d@������������������������       �        �             b@������������������������       �                     4@������������������������       �        ?            �O@'       (                    �?���*ñ?�
           ��@������������������������       �        �
           R�@)       ,                  H�IV@�/����?&             C@*       +                 �56B@�;C�M��?             9@������������������������       �                     7@������������������������       �                      @������������������������       �                     *@�t�b�values�hhK ��h��R�(KK-KK��hX�B�       "�@     ^�@     ƭ@     ؐ@     ܬ@      n@     ��@              ?@      n@      3@              (@      n@      @     �l@             �l@      @              "@      (@              (@      "@             @]@     0�@      Q@      $@      Q@                      $@     �H@     ��@      $@     ��@             ��@      $@             �C@      @     �C@                      @     �e@     �@     �b@      h@      @     �[@       @     @[@             @[@       @              @      �?      @                      �?      b@     �T@      b@      4@      b@                      4@             �O@      7@     p�@             R�@      7@      .@      7@       @      7@                       @              *@�t�bub�_sklearn_version��0.24.2�ub.