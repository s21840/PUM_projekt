���     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �min_impurity_split�N�class_weight�N�	ccp_alpha�G        �_sklearn_version��0.24.2�ub�n_estimators�K
�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�auto�hNhG        hNhG        �n_features_in_�K�n_features_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h-�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh%hNhJ�
hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��h6�f8�����R�(Kh:NNNJ����J����K t�b�C              �?�t�bh>h*�scalar���h9C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hK�
node_count�M�nodes�h,h/K ��h1��R�(KM��h6�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hkh9K ��hlh9K��hmh9K��hnhJK��hohJK ��hph9K(��hqhJK0��uK8KKt�b�BXv         x                  �A��֨4c�?�#         ��A       �                    �?��FK_N�?a�         ��A                           �?���_��?s_          ���@                           �?p��)H�?p!          �i�@                         �HA0�&�ar�?b          ���@������������������������       �        K           ��@       
                   �v�@L��o�?           ��@       	                    �? mčK��?           ��@������������������������       �        �           p�@������������������������       �        E            @Y@������������������������       �                      @                         N�A .���z?           ��@                         `tA ���`;?�           ��@������������������������       �        �           q�@                         �uA����e��?*            �P@������������������������       �                     �?������������������������       �        )            @P@                         �A��ga�=�?(            �P@������������������������       �        !             J@������������������������       �                     .@       V                  xA�豝v�?>          ���@       1                    ��@�a*��?=           (�@                         @"�@���G�?�            �x@                           (p@z�G�z�?             @������������������������       �                     @                           Pu@      �?              @������������������������       �                     �?������������������������       �                     �?       ,                  (�A� �A��?�            Px@       '                  �pA�K1T:�?�            @m@       &                   ��@�����ߒ?z            �j@        %                    �?pY���D�?0            �S@!       $                    �?��?^�k�?+            �Q@"       #                  �LA�nkK�?             G@������������������������       �                     F@������������������������       �                      @������������������������       �                     8@������������������������       �                     "@������������������������       �        J             a@(       +                    8�@�KM�]�?             3@)       *                  �2�@�X�<ݺ?             2@������������������������       �                     �?������������������������       �                     1@������������������������       �                     �?-       0                    �?z�G�z�?^            `c@.       /                  \:A@ެ[�>�?R            @`@������������������������       �        @            �X@������������������������       �                     ?@������������������������       �                     9@2       3                   HA��x�y�?<          ���@������������������������       �        6          �o�@4       7                  ��A4u���?           ��@5       6                    �?p�A�>��?           z@������������������������       �                   �x@������������������������       �                     6@8       M                    �?���H��?�           ؞@9       :                  ��A�F��B��?           X�@������������������������       �                     @;       L                   �A`����E�?           H�@<       =                    �@�r����?�           H�@������������������������       �                     @>       K                   �A�cLN�)�?�           <�@?       H                  �A,0d���?�           8�@@       E                   ��@���:��?           ��@A       D                    ��@�����H�?             "@B       C                   ���@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @F       G                    �?�u����?           ��@������������������������       �        �           ��@������������������������       �        ;            �V@I       J                    �?&P�N�?�            �t@������������������������       �        �            �q@������������������������       �        #             K@������������������������       �                     �?������������������������       �        '             P@N       Q                  �A�H�m�?�            �@O       P                    �?HӘu���?�           H�@������������������������       �        �           0�@������������������������       �        .            �P@R       U                   ��@�LQ�1	�?             7@S       T                    �?���y4F�?
             3@������������������������       �        	             .@������������������������       �                     @������������������������       �                     @W       �                   �L�@h雠�ʽ?�            0y@X       o                    �?�Pk�w��?�             y@Y       ^                  l�A�7��?�            q@Z       ]                  �
A�<ݚ�?             ;@[       \                   ���@      �?
             0@������������������������       �                     @������������������������       �                     $@������������������������       �                     &@_       n                   �{�@`J����?�            �n@`       m                    ��@�YX�Z�?g            �d@a       f                  |�@h㱪��?e            �d@b       e                  �9�@��-�=��?            �C@c       d                    �?�˹�m��?             C@������������������������       �                    �A@������������������������       �                     @������������������������       �                     �?g       h                  p�A ������?J            �_@������������������������       �        =            �Y@i       j                    �@�8��8��?             8@������������������������       �        
             0@k       l                  �A      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �        2            �S@p       s                  ��@��b�h8�?S            �_@q       r                   ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @t       u                  ��@Hn�.P��?Q             _@������������������������       �                    �D@v       �                   Ч�@�+Ĺ+�?8            �T@w       �                  �A ��WV�?5            �S@x       {                    s�@��(\���?             D@y       z                    N�@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @|                         ��A�g�y��?             ?@}       ~                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     9@������������������������       �                     C@�       �                  �A���Q��?             @�       �                  �A�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?ȤP�L��?�         ��A�       �                    �?�1�o�?�         XzA�       �                  �A ��`#g?��          �	�@�       �                  N�A  ��7�?~�           n�@�       �                    �? �����?�          �Z�@�       �                  ԰A  
��?�|          ���@������������������������       �        �{          �|�@�       �                  ��A "���?�            pp@������������������������       �                     �?������������������������       �        �            `p@������������������������       �        �           �@�       �                  p�A@���I�?g            �c@������������������������       �                     �?������������������������       �        f            �c@�       �                  N�A �G�H
�?=           ܴ@������������������������       �                     �?�       �                  $�A�.�����?<           ۴@�       �                  �vA ��w�?�           ̳@������������������������       �        Z           �@�       �                    �?`<)�+�?4            @S@������������������������       �        2            �R@������������������������       �                     @�       �                   ���@�ne�!2�?�            �p@������������������������       �                      @�       �                  �zA`=��?��?�            �p@������������������������       �        �            Pp@������������������������       �                      @�       �                  xA`��&�?P         ���@�       �                  :HAL,��+��?8         P��@������������������������       �        ��          ���@�       �                    �?&�`�.�?�          ���@������������������������       �        �          ���@������������������������       �        �           p�@�       �                    �?�P�<��?           $�@������������������������       �        �           x�@�       �                   �?�@�� ND��?j            `e@������������������������       �                      @�       �                   .�A0u��Fs�?i             e@�       �                  ��A������?E            @[@�       �                   �A�nkK�?              G@�       �                  �(A�C��2(�?             6@������������������������       �                     4@������������������������       �                      @������������������������       �                     8@�       �                   ܻAd�;lr�?%            �O@�       �                  %A�y��*�?"             M@������������������������       �                    �I@������������������������       �                     @�       �                   �Az�G�z�?             @������������������������       �                      @�       �                   �QA�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                  :�A �.�?Ƞ?$             N@������������������������       �        #            �M@������������������������       �                     �?�       �                  6HA��Td��?��           �@������������������������       �        ��          ���@�       u                 ZwA���;+"�?G           "�@�       ,                 \FAJ����8�?�          ���@�       �                   |XA��M�I��?�           ɲ@�       �                  z�A>�Epz�?�	           �@�       �                    �?`x�%�F�?H	           �@������������������������       �                   Ē@�       �                   <�	A��]��/�?<           ��@�       �                    �?�Yr��e�?�           4�@������������������������       �        X           ��@������������������������       �        k            �e@�       �                  �Ax�f� �?y           ��@�       �                   �	A��ػ[�?t           X�@�       �                    �?�+�����?Y           �@������������������������       �        0           ��@������������������������       �        )            �H@�       �                   �A؇���X�?             E@�       �                   �A�q�q�?             @������������������������       �                     �?�       �                   ��@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   6A��-�=��?            �C@������������������������       �        	             0@�       �                    �?�㙢�c�?             7@������������������������       �                     3@������������������������       �                     @�       �                   ��A�q�q�?             @������������������������       �                      @�       �                  �*A      �?             @������������������������       �                      @������������������������       �                      @�       �                  (��@���Q��?Q            @_@�       �                   ��@z�J��?             �G@�       �                    �?h+�v:�?             A@������������������������       �                     5@������������������������       �        
             *@�       �                    �?8�Z$���?
             *@������������������������       �                      @������������������������       �                     &@�       �                  ��A�q�q�?1            �S@�       �                    �?|�U&k�?.            �R@������������������������       �                     G@�       �                   ءA�>4և��?             <@�       �                  �A�q�q�?             (@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                  2�A؇���X�?             @�       �                   Hr�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     0@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       +                   �?d��ȍ�?d           �@�       �                   ��A^���8D�?           ��@�       �                    �?�z�G��?             >@������������������������       �                     5@������������������������       �                     "@�                        |/AB�����?           ��@                         �dAZ4��?�           ��@                         �?��7	C)�?           @z@������������������������       �        u             f@������������������������       �        �            �n@                        �A�d��G��?�            `j@      
                 2�A��"�ű�?�            �i@                       �x�@      �?             6@������������������������       �                     @      	                   �?ҳ�wY;�?             1@������������������������       �                     @������������������������       �                     &@                        �Aܖ�DR�?p            �f@                       ���@>��C��?C             ]@                       ���@^����?1            �U@                        ��A0,Tg��?0             U@                         �?V������?+            �R@������������������������       �                     6@������������������������       �                     J@������������������������       �                     $@������������������������       �                      @                        rA(;L]n�?             >@                       أA      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     <@                         �?�%o��?-            �P@������������������������       �                     5@������������������������       �                      G@                       �Ar�q��?             @������������������������       �                     �?������������������������       �                     @      $                 ��A$Z9��?p            �d@       #                 �qAI����?f            @c@!      "                   �?���3`��?_            �a@������������������������       �                     =@������������������������       �        J             \@������������������������       �                     *@%      &                  J-A�n_Y�K�?
             *@������������������������       �                     @'      *                  dA      �?             $@(      )                 RA      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �        L             `@-      X                  �4ADji3��?�           ��@.      3                 ��A������?�           ��@/      0                   �?�|���v�?           :�@������������������������       �        ;           �@1      2                   �?L�F��?D           ��@������������������������       �        �           ��@������������������������       �        �            0s@4      W                   �?���|���?<             V@5      >                  @&�@�'�=z��?.            �P@6      ;                 *}A �o_��?             9@7      8                 �CA@4և���?             ,@������������������������       �                     "@9      :                   �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?<      =                   �?�eP*L��?             &@������������������������       �                     @������������������������       �                     @?      H                 J�AhP�vCu�?!            �D@@      A                  4A�n_Y�K�?
             *@������������������������       �                     @B      G                  �%Az�G�z�?             $@C      D                  �)A�����H�?             "@������������������������       �                     @E      F                   �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?I      R                 ��A����X�?             <@J      M                 &�A��<b���?             7@K      L                   �?�IєX�?             1@������������������������       �                     �?������������������������       �                     0@N      Q                 P�A�q�q�?             @O      P                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @S      T                  �^A���Q��?             @������������������������       �                     �?U      V                 ��A      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     6@Y      p                  h�Af�Sc��?;            �X@Z      _                  �BA����X�?3             U@[      \                 B�A�}�+r��?             3@������������������������       �                     .@]      ^                   �?      �?             @������������������������       �                     @������������������������       �                     �?`      a                   �?�y(dD�?-            @P@������������������������       �                    �@@b      i                  n^A     ��?             @@c      h                  �VA      �?             0@d      e                 Ġ	A"pc�
�?	             &@������������������������       �                     �?f      g                   �?ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     @j      m                 �A     ��?             0@k      l                   �?      �?              @������������������������       �                      @������������������������       �                     @n      o                   �?      �?              @������������������������       �                     @������������������������       �                     �?q      r                  ^�A؇���X�?             ,@������������������������       �                     @s      t                  ԓA����X�?             @������������������������       �                      @������������������������       �                     @v      w                   �?�����H�?T            �`@������������������������       �        K             ^@������������������������       �        	             .@y                         �?�A���?](          ���@z      �                  
`A�Pq����?I           ��@{      �                   �?��Z@t�?�           ��@|      �                 }A�G60��?�           6�@}      ~                 pGAd㯅��?�           �@������������������������       �        	           ��@      �                   �?cde�?�            p@������������������������       �        �            `l@������������������������       �                     >@�      �                   �?��hJ,�?             A@������������������������       �                     =@������������������������       �                     @�      �                 j#AxUV�	��?           ��@�      �                  �Ah���*C�?=	           &�@������������������������       �        9             X@�      �                 $�A0��<��?	           f�@�      �                 ���@� .&8>�?�           ��@�      �                 �A���E0�?�           P�@�      �                 ���@�2s��?�           8�@�      �                 г�@�Q����?�           (�@�      �                 (^�@�]0��<�?K            �^@�      �                  �@�ȉo(��?>            �V@�      �                  ��@(;L]n�?=            �V@�      �                   �?P�2E��?.            @P@������������������������       �        +             O@������������������������       �                     @������������������������       �                     9@������������������������       �                     �?������������������������       �                     ?@�      �                 ��@<J96���?�           X�@�      �                   �? ���g=�?�           h�@������������������������       �        _           (�@������������������������       �        *             R@�      �                 ��@�z�G��?             >@������������������������       �                     @�      �                  ,�A�J�4�?             9@�      �                  :�A�q�q�?             @������������������������       �                      @�      �                 (2�@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     3@������������������������       �                      @������������������������       �                     @�      �                 �A���ّ��?�           ܖ@�      �                 �1A�2��Ǫ�?�           Ė@�      �                   �?`�}�O�?@           0�@������������������������       �                   ��@������������������������       �        $            �I@�      �                 �<A(L�\�?j           X�@������������������������       �                     @�      �                 ܁A0�<jX��?i           8�@�      �                 ,tA��T\��?�            �s@�      �                 t%
AD�/�6��?�            �s@�      �                  ̛A��`T.1�?�            �k@������������������������       �                     �?�      �                   �?t��ճC�?�            �k@������������������������       �        �            �i@������������������������       �        
             .@�      �                   �?��k=.��?@            �W@������������������������       �        5             S@������������������������       �                     2@������������������������       �                      @�      �                 8OA0��d��?�            @m@������������������������       �        '             O@�      �                   �?�Ts�k��?p            �e@������������������������       �        i             d@������������������������       �                     &@�      �                   �?�q�q�?             @������������������������       �                     @������������������������       �                      @�      �                  ΝA,�Y���?m           ȕ@�      �                 ��AX�Cc�?	             ,@�      �                 ���@�q�q�?             @������������������������       �                      @������������������������       �                     @�      �                   �?      �?              @������������������������       �                     @������������������������       �                     �?�      �                   �? ���g=�?d           ��@������������������������       �                   �@������������������������       �        b             d@�      �                 @�AP&��H��?�           ��@�      �                 x�@@c����?�            @u@������������������������       �        t             g@�      �                 �0�@�(�Tw�?b            �c@������������������������       �                     �?�      �                 ��A u�z\A�?a            `c@������������������������       �        /            �S@�      �                   �?�"w����?2             S@������������������������       �        .             R@�      �                 DA      �?             @������������������������       �                     �?������������������������       �                     @�      �                 fBA Os���?�             z@�      �                 �;A�8��?f            �d@�      �                   �?�nkK�?a             d@������������������������       �        Z            @c@������������������������       �                     @�      �                   �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        �            `o@�                         �?�(����?�	           �@�      �                 �xA5$'{�?r           �@�      �                 `��@��Q�w��?d           ��@�      �                  ��A���*~�?:            @V@�      �                 �A�+$�jP�?4            @T@������������������������       �        +            @P@�      �                   �?      �?	             0@������������������������       �                     .@������������������������       �                     �?�      �                 (+A      �?              @������������������������       �                     @������������������������       �                     @�      �                  ��A�?�N
�?*           \�@�      �                 %�@�6����?'           D�@�      �                 �@A�R��#�?�            �i@������������������������       �        }            @i@������������������������       �                     @�      �                 BMA��g�?�           �@������������������������       �        q           x�@�      �                  f�A�5U��K�?4            �T@������������������������       �        $            �L@�      �                 [�@�	j*D�?             :@������������������������       �                      @�      �                   �?      �?             8@������������������������       �        
             2@������������������������       �                     @�      �                 ��A�q�q�?             @������������������������       �                     @������������������������       �                      @�      �                  ̳A���7�?             6@������������������������       �                     .@�                          �?؇���X�?             @������������������������       �                     @������������������������       �                     �?                         �?P����>�?           �@������������������������       �        b           �@                       VIA �Zz�q�?�            �p@������������������������       �        �            @m@������������������������       �                     ?@                       yA(��n�?           �@                         �?�	��ϋ�?�           ��@	                         �@�~Zd��?           ��@
                        r�A������?D             [@                        ,vA�ջ����?A             Z@������������������������       �        1            @T@                         �?�nkK�?             7@������������������������       �                     $@                        ��@$�q-�?
             *@������������������������       �                     @                        �Ar�q��?             @������������������������       �                     �?������������������������       �                     @                        �A      �?             @������������������������       �                      @������������������������       �                      @                       zFA({���?;           6�@������������������������       �        
           O�@������������������������       �        1           p~@������������������������       �        ]           ��@                         �? �\���?8            �S@������������������������       �        4            �R@������������������������       �                     @�t�b�values�h,h/K ��h1��R�(KMKK��hJ�B�!      �!A    ���@    |�A    ���@    @D�@     ȩ@    ���@     ��@     �@     p�@     ��@             �Y@     p�@     @Y@     p�@             p�@     @Y@               @             �@      0@     ��@      �?     q�@             @P@      �?              �?     @P@              J@      .@      J@                      .@    @�@     �@     �@     �@     @u@      K@      �?      @              @      �?      �?      �?                      �?     0u@      I@     �j@      3@     �j@       @     @S@       @      Q@       @      F@       @      F@                       @      8@              "@              a@               @      1@      �?      1@      �?                      1@      �?              _@      ?@     �X@      ?@     �X@                      ?@      9@             ��@     ��@    �o�@             p@     ��@      6@     �x@             �x@      6@             `m@     ,�@      d@     ؐ@      @             �c@     ؐ@     �c@     ��@      @              c@     ��@      c@     ��@     �X@     �@       @      �?       @      �?       @                      �?      @             �V@     ��@             ��@     �V@              K@     �q@             �q@      K@              �?                      P@     �R@     ��@     �P@     0�@             0�@     �P@               @      .@      @      .@              .@      @              @              9@     �w@      6@     �w@      ,@     0p@      @      5@      @      $@      @                      $@              &@       @     �m@       @     �c@      @     �c@      @     �A@      @     �A@             �A@      @              �?               @      _@             �Y@       @      6@              0@       @      @       @                      @       @                     �S@       @     �]@       @      �?              �?       @              @     �]@             �D@      @     @S@      @     �R@      @     �B@       @      @              @       @              �?      >@      �?      @              @      �?                      9@              C@      @       @      �?       @      �?                       @       @              @            ��A    �k�@    (�A     ��@    ���@     �U@    �m�@       @    `Z�@      �?    ���@      �?    �|�@             `p@      �?              �?     `p@             �@             �c@      �?              �?     �c@             ��@     @U@              �?     ��@      U@     ��@     �R@     �@              @     �R@             �R@      @             Pp@      $@               @     Pp@       @     Pp@                       @    ���@    ���@    @��@    ���@    ���@             p�@    ���@            ���@     p�@             `c@     ��@             x�@     `c@      0@               @     `c@      ,@      X@      *@      F@       @      4@       @      4@                       @      8@              J@      &@     �I@      @     �I@                      @      �?      @               @      �?       @      �?                       @     �M@      �?     �M@                      �?    ���@     H�@    ���@             ��@     H�@     گ@     е@      �@     ��@     ��@     T�@     \�@     �@     Ē@             �l@     �@     �e@     ��@             ��@     �e@             �L@     ��@     �K@     ��@     �H@     ��@             ��@     �H@              @      B@       @      �?      �?              �?      �?      �?                      �?      @     �A@              0@      @      3@              3@      @               @      @               @       @       @       @                       @     �R@      I@      7@      8@      5@      *@      5@                      *@       @      &@       @                      &@      J@      :@     �I@      7@      G@              @      7@      @      @      @      �?              �?      @              �?      @      �?       @               @      �?                      @              0@      �?      @      �?                      @     `z@     ��@     Pr@     ��@      5@      "@      5@                      "@      q@     p�@     �m@     �x@      f@     �n@      f@                     �n@      O@     �b@     �L@     �b@      &@      &@      @              @      &@      @                      &@      G@      a@      9@     �V@      8@      O@      6@      O@      6@      J@      6@                      J@              $@       @              �?      =@      �?      �?              �?      �?                      <@      5@      G@      5@                      G@      @      �?              �?      @              A@     �`@      =@     @_@      =@      \@      =@                      \@              *@      @       @              @      @      @      @      @              @      @                       @      `@             ʠ@     �@     N�@     ֤@     ��@     ��@     �@             0s@     ��@             ��@     0s@              L@      @@      A@      @@      2@      @      *@      �?      "@              @      �?      @                      �?      @      @      @                      @      0@      9@       @      @              @       @       @       @      �?      @              @      �?      @                      �?              �?       @      4@      @      2@      �?      0@      �?                      0@      @       @      �?       @      �?                       @      @              @       @              �?      @      �?              �?      @              6@              O@      B@      N@      8@      2@      �?      .@              @      �?      @                      �?      E@      7@     �@@              "@      7@       @      ,@       @      "@      �?              �?      "@              "@      �?                      @      @      "@      @       @               @      @              �?      @              @      �?               @      (@              @       @      @       @                      @      .@      ^@              ^@      .@             ��@     ]�@     �@     (�@      �@     �@     6�@      p@     ,�@     `l@     ��@              >@     `l@             `l@      >@              @      =@              =@      @             Pw@     �@     pv@     X�@              X@     pv@     ��@     @h@     ��@     �V@     ��@     �U@     ��@     @U@     ��@      @     �]@      @     �U@      @     �U@      @      O@              O@      @                      9@      �?                      ?@     @T@     Ё@      R@     (�@             (�@      R@              "@      5@      @              @      5@      @       @       @               @       @       @                       @              3@       @              @              Z@     <�@     �Y@     ,�@     �I@     ��@             ��@     �I@             �I@     �@      @             �G@     �@      B@     �q@      A@     �q@      0@     �i@      �?              .@     �i@             �i@      .@              2@      S@              S@      2@               @              &@     �k@              O@      &@      d@              d@      &@               @      @              @       @             �d@     4�@      @      "@      @       @               @      @              �?      @              @      �?              d@     �@             �@      d@              ,@     @�@       @      u@              g@       @     @c@      �?              �?     @c@             �S@      �?     �R@              R@      �?      @      �?                      @      (@     `y@      (@     `c@      @     @c@             @c@      @              @      �?              �?      @                     `o@     З@     (�@     (�@      _@     $�@     �Y@     �Q@      3@     �P@      .@     @P@              �?      .@              .@      �?              @      @      @                      @     �@      U@     �@      T@     @i@      @     @i@                      @     ��@     �R@     x�@               @     �R@             �L@       @      2@       @              @      2@              2@      @               @      @              @       @              �?      5@              .@      �?      @              @      �?             @m@     0�@             �@     @m@      ?@     @m@                      ?@     ڳ@     ��@     ֳ@     �~@     ��@     �~@     @Z@      @     �Y@      �?     @T@              6@      �?      $@              (@      �?      @              @      �?              �?      @               @       @               @       @             O�@     p~@     O�@                     p~@     ��@              @     �R@             �R@      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ/��hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaM�hbh,h/K ��h1��R�(KM���hi�B�]         �                  BHA�C��?�#         ��A       ?                    �?�vZ���?��         p�A                           �?`��8���?�U          `��@������������������������       �                  ���@       6                  �6A@�`s�@�?�7           ��@                         xA�޲��r�?'0          ���@������������������������       �        e/          ���@       /                    �?0����a�?�            �s@	                         ���@��JB��?�            �i@
                         ���@���Q��?             $@������������������������       �                     @������������������������       �                     @                         <�APKvke�?            �h@                           �?�q�q�?             5@������������������������       �        
             ,@������������������������       �                     @       ,                  ��A����k��?q             f@                         ���@86��Z�?e            �c@������������������������       �                     :@       %                   �S�@�U�=���?U            �`@                         ���@`Jj��?O             _@������������������������       �                     �?       "                  ��@��sK�z�?N            �^@                          ���@؇���X�?            �A@                         d�A�q�q�?             (@                         ���@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @       !                  p��@�nkK�?             7@                            ��@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             1@#       $                    �?`���i��?<             V@������������������������       �        :            �U@������������������������       �                      @&       '                   �h�@      �?              @������������������������       �                     �?(       )                    J�@؇���X�?             @������������������������       �                     @*       +                  �A�q�q�?             @������������������������       �                     �?������������������������       �                      @-       .                    �?�E��ӭ�?             2@������������������������       �        	             *@������������������������       �                     @0       3                    ��@(N:!���?>            @Z@1       2                    �?      �?             @������������������������       �                     �?������������������������       �                     @4       5                    �?��T�u��?<            @Y@������������������������       �        5             W@������������������������       �                     "@7       8                  $wA�\K��?v           ��@������������������������       �        Q           �@9       :                    \�@���7�?%            �P@������������������������       �                      @;       <                    �?     ��?$             P@������������������������       �                     H@=       >                  (�A      �?             0@������������������������       �        
             .@������������������������       �                     �?@       �                   &�A������?�z         �lAA       |                   �1A���n���?�V         �AB       {                    �?�ft�?�         ��AC       D                    �? Ja7��?��          ���@������������������������       �        �V          �>�@E       b                  N�A��cB���?�          P�@F       O                  txA�k^|�?+�          `��@G       N                    �? @�4�3?6�          � �@H       M                  ���@ @8��P?j          �3�@I       J                   �
A h���a0?P'          �@�@������������������������       �        �           ?�@K       L                   <�
A ���BR?�           �@������������������������       �                      @������������������������       �        �           �@������������������������       �        X          `c�@������������������������       �        �           h�@P       S                  &�A�2s��?�           8�@Q       R                    �?`�рv�?�           0�@������������������������       �        �           �@������������������������       �        )            @Q@T       _                  ̕A
��[��?+            @P@U       Z                   lIA      �?
             0@V       W                  ƺAףp=
�?             $@������������������������       �                     @X       Y                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @[       \                   �
Ar�q��?             @������������������������       �                     @]       ^                  >A      �?              @������������������������       �                     �?������������������������       �                     �?`       a                    �?ZՏ�m|�?!            �H@������������������������       �                    �D@������������������������       �                      @c       t                   ��@`�Gc�?�           Z�@d       e                  �wA�H�I���?           l�@������������������������       �        �           2�@f       o                  ��A>���Rp�?             =@g       h                  ��A��2(&�?             6@������������������������       �                     $@i       j                    ��@      �?             (@������������������������       �                     �?k       l                  ʯA"pc�
�?             &@������������������������       �                     @m       n                    �?      �?             @������������������������       �                      @������������������������       �                      @p       s                  �Aև���X�?             @q       r                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @u       v                   ��@p2'*�?�           ��@������������������������       �                      @w       z                    �?��u���?�           ��@x       y                  6vA01-�W��?�
           а@������������������������       �        \
           |�@������������������������       �        2             U@������������������������       �        $            }@������������������������       �        ӆ          @��@}       ~                   �1A �Hd�e�?��           I�@������������������������       �                     @       �                    �? j��B�?��          �H�@�       �                  LxA��@c&��?��          �n�@������������������������       �        [�          ���@�       �                  |]A���� �?K           �@�       �                    �?j����?�           ��@�       �                   ��A������?�           ��@�       �                   LA9v#4^�?a           ��@�       �                    �?f�t����?�             q@������������������������       �        C            �Z@������������������������       �        l            �d@�       �                   �#A$⍮�l�?�            r@�       �                   �nA��%��?�            �i@�       �                    �?6�iL�?N            �]@������������������������       �                     @@������������������������       �        9            �U@�       �                  ��@��T|n�?2            �U@�       �                    �?�q�q�?
             (@������������������������       �                     @������������������������       �                     @�       �                    �?������?(            �R@������������������������       �                      @������������������������       �        %            �P@�       �                  *|A������?2            @U@������������������������       �                     @�       �                    �?���Q��?0             T@������������������������       �                     @@������������������������       �                      H@�       �                    �?�~����?V            �`@������������������������       �        '            @P@������������������������       �        /             Q@������������������������       �        >             X@�       �                   N�A:wXFpw�?V            �`@�       �                    �?L� P?)�?>            @X@������������������������       �                     1@�       �                    �?�(\����?3             T@������������������������       �        1            �S@������������������������       �                      @�       �                  n�A�\��N��?             C@�       �                   D!Ar�q��?             2@�       �                  ��A      �?             @������������������������       �                     @������������������������       �                     @������������������������       �        	             (@�       �                    �?R���Q�?             4@������������������������       �                     @������������������������       �        	             1@������������������������       �        &L          @F�@�       �                    �?&`�ւ�?z$           ��@�       �                    �?`���/�?t           ��@�       �                  &A����٘?0           }�@�       �                  �xA�h%�M��?           ^�@������������������������       �        �
           *�@������������������������       �        "             J@�       �                  N'A��a�n`�?             ?@������������������������       �                     �?�       �                    �?��S�ۿ?             >@������������������������       �                     5@�       �                  �8A�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �        D           �@�       �                    �?��Xj�?           �@�       �                  &�A �(���?�           ��@�       �                  ��A|~%+�O�?�           �@�       �                   bdA�v�?�?�           �@�       �                    �?|���J��?l	           ҭ@������������������������       �        �           �@������������������������       �        �            0v@�       �                    �?���4�?           2�@������������������������       �        �           ��@������������������������       �        �             n@������������������������       �                      @�       �                    �?��§�ͺ?           �y@������������������������       �        �            �x@������������������������       �                     7@�       �                  �BA�����?w           �@�       �                   `#A@$�.�l�?           �@�       �                  ���@`��* *�?�           (�@������������������������       �        �            �w@�       �                   ޶A��̍$��?�           <�@�       �                    �?�w���l�?�            Pp@�       �                  ��@ :��?�            �l@������������������������       �                     @�       �                   ,�AЇ�γ��?�            �l@�       �                  (yA@3�qH�?h             d@������������������������       �        I            �\@�       �                  �EA��<b�ƥ?             G@������������������������       �                    �F@������������������������       �                     �?�       �                  �qA�L#���?.            �P@������������������������       �        ,            �O@������������������������       �                     @������������������������       �                     >@�       �                    �?��.���?
           P�@�       �                  0wA� ��I�?�           ��@������������������������       �        �           p�@������������������������       �                     @������������������������       �        '             K@�       �                   �#A �-�_��?~           ��@������������������������       �                      @�       �                  �zA��,�b��?}           ��@������������������������       �        m           �@�       �                  J�A�X�<ݺ?             B@������������������������       �                     >@�       �                  ��A�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   �dA@4և���?a            @c@�       �                   ��A@�E�x�??            �X@�       �                   ��A���7�?             6@������������������������       �                     5@������������������������       �                     �?�       �                    �?�"w����?1             S@�       �                  �CA`����֜?,            �Q@������������������������       �                     �?������������������������       �        +            @Q@������������������������       �                     @�       �                   �gA�X�C�?"             L@������������������������       �                     @�       �                    �?���C��?!            �J@�       �                  r�A�t����?            �I@������������������������       �                    �F@������������������������       �                     @������������������������       �                      @�       h                   �?j+���?�R           R�@�                          �?>v��??J          @<�@�                          �?�= ���?�           ^�@�       �                    �?Dp'r��?�           ��@������������������������       �        �           ��@                         �G�@ R�,3��?           �y@������������������������       �        T            �^@                        ���@��VYw��?�            �q@������������������������       �                      @      	                 �pA r���?�            �q@                       *nA��<�Ұ?a            `b@                       :^A�k~X��?`             b@������������������������       �        _            �a@������������������������       �                      @������������������������       �                     @
                       �YA�Ŗ�Pw�?Z            @a@������������������������       �        Y             a@������������������������       �                     �?������������������������       �        �           �@      9                 `A�,ٱ-��?�A          ���@      8                   �?���K�E�?x            �@                       �HA�m�Hɷ?�            Px@                       �|�@      �?              @������������������������       �                     @                       ~HAz�G�z�?             @                       NHA      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @      7                 �wA�m(']�?�            �w@                         �@�UM���?�            �w@                       �\A�θ�?             *@                        [�@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?                       ^A�q�q�?             @������������������������       �                      @������������������������       �                     �?!      "                 �OAp��ӵ6�?�            �v@������������������������       �        <             Z@#      2                   �?؀���˲?�            `p@$      %                 �OAXpBt,��?t            �e@������������������������       �                     �?&      +                 \CA`��F:u�?s            �e@'      *                 4;ADu9iH��?8            �U@(      )                  �CA���N8�?7             U@������������������������       �        4             T@������������������������       �                     @������������������������       �                      @,      -                 `[A`���i��?;             V@������������������������       �        (             O@.      /                 d�A$�q-�?             :@������������������������       �                     0@0      1                  |�Az�G�z�?             $@������������������������       �                      @������������������������       �                      @3      6                 DSA���E�?5            �U@4      5                 �RA@4և���?
             ,@������������������������       �        	             *@������������������������       �                     �?������������������������       �        +            @R@������������������������       �                      @������������������������       �        �           ��@:      g                   �?r�'����?'?          ���@;      f                 �xA�[貎�?�           �@<      _                 :gA����y��?�          ���@=      T                   �?��� *�?o           ��@>      O                 ��AتNq
�?j	           ĭ@?      L                 ĕA�o����?f	           ��@@      C                  {@�U��^�?l           ��@A      B                 �UA      �?             @������������������������       �                      @������������������������       �                      @D      G                 H�AȋJ�0B�?j           ��@E      F                  V�A 8b.���?,           ��@������������������������       �        �           �@������������������������       �        �             k@H      I                 ��A ���x�?>            @\@������������������������       �                      @J      K                  �A��E�wx�?=            �[@������������������������       �        7            �X@������������������������       �                     *@M      N                  0�ApY���D�?�            �x@������������������������       �        �            x@������������������������       �                     $@P      S                 @�Aև���X�?             @Q      R                  D�Az�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @U      X                 �aA�2�~w�?           �@V      W                 �`A���Q��?             @������������������������       �                      @������������������������       �                     @Y      \                 �UA�6�ػ?           ܞ@Z      [                  �Ap�]�&9�?            Ȟ@������������������������       �        �           �@������������������������       �        J            �[@]      ^                 �A���Q��?             @������������������������       �                     @������������������������       �                      @`      c                   �?�<'L���?&           2�@a      b                  ��A=�F	��?w           ��@������������������������       �        J           ��@������������������������       �        -            �O@d      e                  ��A �#�Ѵ�?�           ̐@������������������������       �        �           �@������������������������       �        %             I@������������������������       �        J            �[@������������������������       �        H)           V�@i      �                 �}A`��PE?�?�           >�@j      o                  z�A��S^��?�           �@k      l                   �? �����C?"           ĩ@������������������������       �        �           ��@m      n                 lvA �o�8O?5           d�@������������������������       �        4           b�@������������������������       �                     �?p      }                 ��A��q���?_            �a@q      r                   �?�f7�z�?;            �U@������������������������       �                     E@s      z                 �Az�G�z�?             �F@t      w                 
iA��-�=��?            �C@u      v                   �?�IєX�?             A@������������������������       �                     @@������������������������       �                      @x      y                   �?���Q��?             @������������������������       �                     @������������������������       �                      @{      |                   �?r�q��?             @������������������������       �                     �?������������������������       �                     @~      �                 X]A      �?$             L@      �                 ,vA��a�n`�?             ?@�      �                  ƛA���Q��?             $@�      �                   �?և���X�?             @�      �                 ��A      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�      �                  v�A؇���X�?             5@������������������������       �                     �?�      �                   �?ףp=
�?             4@������������������������       �                     �?�      �                 �A�}�+r��?             3@�      �                  �Az�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     ,@�      �                 A� �	��?             9@�      �                 �A
;&����?             7@�      �                   �?ҳ�wY;�?
             1@������������������������       �                     @�      �                  DA��
ц��?             *@�      �                   �?����X�?             @������������������������       �                     @������������������������       �                      @�      �                   �?r�q��?             @������������������������       �                     �?������������������������       �                     @�      �                   �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�      �                 b�A��c:�?             G@�      �                   �?p9W��S�?             C@�      �                   �?$�q-�?             :@������������������������       �                     @�      �                 \�A�C��2(�?             6@�      �                 ʗA���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     1@�      �                   �?      �?             (@������������������������       �                      @�      �                 T�Aףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                      @�t�bh~h,h/K ��h1��R�(KM�KK��hJ�B�      �A     ��@    �^A     :�@    @��@     u@    ���@            ���@     u@    @��@      q@    ���@              C@      q@      :@     �f@      @      @              @      @              6@     �e@      @      ,@              ,@      @              .@      d@      $@     �b@              :@      $@     �^@       @      ]@      �?              @      ]@      @      >@      @       @      @       @               @      @                      @      �?      6@      �?      @      �?                      @              1@       @     �U@             �U@       @               @      @      �?              �?      @              @      �?       @      �?                       @      @      *@              *@      @              (@     @W@      @      �?              �?      @              "@      W@              W@      "@             $�@     �O@     �@              @     �O@       @              �?     �O@              H@      �?      .@              .@      �?            @�A     �@    (tA     ��@    ��A     ��@    �s�@     ��@    �>�@            ��@     ��@     +�@     ��@    @ �@       @    @3�@       @    �?�@       @     ?�@             �@       @               @     �@            `c�@             h�@             �U@     ��@     @Q@     �@             �@     @Q@              2@     �G@      $@      @      "@      �?      @              @      �?              �?      @              �?      @              @      �?      �?              �?      �?               @     �D@             �D@       @             �@      [@     @�@      6@     2�@              @      6@      @      3@              $@      @      "@      �?               @      "@              @       @       @               @       @              @      @      @      �?              �?      @                       @     N�@     �U@               @     N�@      U@     |�@      U@     |�@                      U@      }@            @��@             '�@      �@              @     '�@     �@    �*�@     �@    ���@              x@     �@     �u@     �{@     `o@     �{@     @g@     pw@     �Z@     �d@     �Z@                     �d@     �S@     @j@     �G@     �c@      @@     �U@      @@                     �U@      .@     �Q@      @      @      @                      @       @     �P@       @                     �P@      @@     �J@              @      @@      H@      @@                      H@     @P@      Q@     @P@                      Q@      X@             �B@     �X@      3@     �S@      1@               @     �S@             �S@       @              2@      4@      .@      @      @      @      @                      @      (@              @      1@      @                      1@    @F�@            ���@     ��@     g�@     �K@     F�@     �K@     *�@      J@     *�@                      J@      <@      @              �?      <@       @      5@              @       @      @                       @     �@             x�@     t�@     `�@     7�@     ��@     ��@     ��@     ��@     0v@     �@             �@     0v@              n@     ��@             ��@      n@               @              7@     �x@             �x@      7@             ��@     �N@     ��@      I@     �@      ,@     �w@             �@      ,@     �o@       @     �k@       @              @     �k@      @      d@      �?     �\@             �F@      �?     �F@                      �?     �O@      @     �O@                      @      >@              �@      @     p�@      @     p�@                      @      K@             �@      B@               @     �@      A@     �@               @      A@              >@       @      @       @                      @     �a@      &@      X@       @      5@      �?      5@                      �?     �R@      �?     @Q@      �?              �?     @Q@              @             �G@      "@              @     �G@      @     �F@      @     �F@                      @       @             �@    ���@     o�@    ���@      y@     :�@      y@     ؈@             ��@      y@       @     �^@             pq@       @               @     pq@      @     �a@      @     �a@       @     �a@                       @              @      a@      �?      a@                      �?             �@     ��@    �}�@      w@     ��@      w@      3@      @      @              @      @      �?      �?      �?      �?                      �?      @             �v@      .@     �v@      *@      $@      @      "@      �?      "@                      �?      �?       @               @      �?             @v@      $@      Z@             �o@      $@     �d@      "@              �?     �d@       @      T@      @      T@      @      T@                      @               @     �U@       @      O@              8@       @      0@               @       @       @                       @     �U@      �?      *@      �?      *@                      �?     @R@                       @             ��@     ڿ@     ��@     ڿ@     `�@     ڿ@     �}@     2�@     �v@     ֫@     �n@     Ϋ@     �n@     ̨@     @m@       @       @               @       @             Ȩ@      m@     �@      k@     �@                      k@     �X@      .@               @     �X@      *@     �X@                      *@     x@      $@     x@                      $@      @      @      @      �?      @                      �?               @     �@     @]@       @      @       @                      @     �@     �\@     �@     �[@     �@                     �[@       @      @              @       @             P�@     @\@     ��@     �O@     ��@                     �O@     �@      I@     �@                      I@             �[@             V�@     x�@     �X@     R�@      R@     ©@      �?     ��@             b�@      �?     b�@                      �?      R@     �Q@     �I@      B@      E@              "@      B@      @     �A@       @      @@              @@       @               @      @              @       @              @      �?              �?      @              5@     �A@      @      8@      @      @      @      @      �?      @      �?                      @      @                      @      @      2@      �?               @      2@      �?              �?      2@      �?      @              @      �?                      ,@      ,@      &@      (@      &@      &@      @      @              @      @       @      @              @       @              @      �?              �?      @              �?      @      �?                      @       @              3@      ;@      &@      ;@       @      8@              @       @      4@       @      @              @       @                      1@      "@      @               @      "@      �?      "@                      �?       @        �t�bub��I     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJu�7hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaM�hbh,h/K ��h1��R�(KM���hi�B�U         d                    �?�!+Up�?�#         ��A       -                    �?@�x��t�?�         ��@                          ,�@�Ȫ���?.!           ��@       	                    y�@�ӭ�a��?-             R@                           �?�q�q�?             "@                         \�A      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     �?
                           �?�[|x��?(            �O@                          �2�@      �?             D@                         BA�8��8��?             B@������������������������       �                    �@@������������������������       �                     @                         *�A      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     7@       ,                    �?XmF��f�?!           ��@                         6IAp��R�U�?�           C�@������������������������       �        �           ��@                         ��A�q4��?�           x�@                           �?�Z���?e           x�@������������������������       �        �            �v@                         �zA�h,mṡ?�            `l@������������������������       �        �            �k@������������������������       �                     @                          �@�8x#��?{           x�@������������������������       �                     @       #                   ���@�(�.Y��?z           `�@       "                   ���@�I��7u�?�            0p@        !                    �?����?�            �o@������������������������       �        e            �d@������������������������       �        ?            @V@������������������������       �                     @$       %                  P,�@N��-%�?�            �t@������������������������       �                     7@&       )                  ��A�ɟ=M�?�             s@'       (                    �?      �?�            @r@������������������������       �        �            `k@������������������������       �        :            @R@*       +                    �?����X�?	             ,@������������������������       �                     @������������������������       �                     $@������������������������       �        =           ��@.       ?                  BHA����{�?p�          �s�@/       0                  �yA �"�,�_?��          ���@������������������������       �        ��          ���@1       2                   v�A0a����?           4�@������������������������       �        �           Ē@3       >                    �?��	,UP�?3             W@4       5                  8lA$�q-�?"            @P@������������������������       �                    �F@6       7                  A      �?             4@������������������������       �                      @8       ;                   ��Ar�q��?             2@9       :                  � A      �?             @������������������������       �                      @������������������������       �                      @<       =                    �?@4և���?             ,@������������������������       �                     *@������������������������       �                     �?������������������������       �                     ;@@       Y                  �xA��VG��?�          �8�@A       X                    �?0n�6Ǹ?c          ���@B       M                  �2APvX0|��?�           ��@C       J                    �?��И��?�           $�@D       G                  2�A�8���?B           ش@E       F                   ��Ah]X����?>           Ӵ@������������������������       �        �           ��@������������������������       �        �             q@H       I                   @�A���Q��?             @������������������������       �                     @������������������������       �                      @K       L                   �A��00`��?S           �@������������������������       �        �           ��@������������������������       �        k            �d@N       W                  ��A��P���?&            �@O       P                  �4A`����U�?%           ��@������������������������       �                     @Q       T                    �?��钲��?$           ؊@R       S                   $�A��;�ڒ�?J           p�@������������������������       �        6           p~@������������������������       �                    �C@U       V                   r�A̹�"���?�            �t@������������������������       �        �            �r@������������������������       �                    �@@������������������������       �                      @������������������������       �        �           ��@Z       a                    �?$�q-�?e            �c@[       ^                  ��A�C��2(�?D            �X@\       ]                    �?Pq�����?<            @U@������������������������       �        :            @T@������������������������       �                     @_       `                    �?X�Cc�?             ,@������������������������       �                     "@������������������������       �                     @b       c                    �?�}�+r��?!            �L@������������������������       �                     K@������������������������       �                     @e       L                   �?pִ�d�??         ��	Af       �                   �A�O����?��         pFAg       �                    �?t
9	�T�?�         hAh       �                    ��@@'�y��?47           ��@i       t                    �?��n�?�            pw@j       s                  A4C��J�?�             n@k       n                  � A�K7_�?�            `i@l       m                  ��A�6H�Z�?I            @]@������������������������       �        H             ]@������������������������       �                     �?o       p                  ԝA���1j	�?8            �U@������������������������       �                     �?q       r                  �APq�����?7            @U@������������������������       �        4            @T@������������������������       �                     @������������������������       �                     C@u       x                    �w@�'݊U�?Q            �`@v       w                  lA�BE����?'             O@������������������������       �                    �D@������������������������       �        
             5@y       �                  .A�n���?*             R@z       �                     �@hA� �?(            �Q@{       |                     �@Pa�	�?%            �P@������������������������       �                    �D@}       ~                  �AHP�s��?             9@������������������������       �                     *@       �                    ă@r�q��?             (@������������������������       �                      @������������������������       �                     $@�       �                  @�A      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    ��@@ҳ�h��?L6          @g�@�       �                  ||A�T|�T��?S           ��@�       �                   @�@��Z�?           ��@�       �                   ��@|T(W�j�?�           ��@�       �                  JJA D�^X�?�           ��@������������������������       �        e           �@������������������������       �        4           �~@������������������������       �                      @�       �                   ���@H�]t��?{           J�@�       �                  \A�X��C�?�            �v@������������������������       �        �            �u@������������������������       �                     3@�       �                    �?��W8 �?�           ��@�       �                    8�@�6v��u�?           D�@�       �                  z�A��مD�?3            @S@�       �                  4�Af.i��n�?            �F@������������������������       �                     ?@������������������������       �                     ,@�       �                  �A     ��?             @@������������������������       �                     =@������������������������       �                     @�       �                   ���@d	��ܐ�?�           �@������������������������       �                    �J@�       �                  �<A�X?%�`�?�           <�@������������������������       �        }           ��@������������������������       �        9            �V@�       �                   @?�@<I����?�           8�@�       �                  :)A �ղ?s            �f@������������������������       �        n             f@������������������������       �                     @�       �                   �H�@��s���?            {@������������������������       �                      @�       �                   @^�@�E����?           �z@�       �                  |KA�%���W�?           @y@������������������������       �        �            �v@������������������������       �                    �D@������������������������       �                     :@������������������������       �        >            �U@�       �                  BHAl�����?�#          �S�@�       �                  �wA@�n�1�?1            d�@������������������������       �        �           ��@������������������������       �        �             j@������������������������       �        �           |�@�       �                  �wA�p�B�?��         �]A�       �                  :HA\���9��?/�         0A������������������������       �        wY         � A������������������������       �        �'          �j�@�       �                    �?D3�f�"�?�           ��@������������������������       �        �           ��@�       �                   P�A|y����?�           @�@�       �                   �A�� =�	�?)            @�       �                  ��A$e���?(           �~@�       �                  �0ANKF����?9            @V@������������������������       �        0             R@������������������������       �        	             1@�       �                   dIA,��]L�?�            @y@�       �                   t7A�ˠ�?�             v@�       �                  ��Aףp=
�?�            �u@�       �                   �x	A���d�?�            �u@�       �                  �gA��T����?�            �s@������������������������       �        �            �q@������������������������       �                     9@�       �                  \kA������?             A@������������������������       �                     :@������������������������       �                      @�       �                  �]A      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     J@������������������������       �                     @�       �                   �A@��z��?�            �s@�       �                   |=ApNho&,�?�            �n@�       �                  ~�A�L��ȕ?C            @W@������������������������       �        B             W@������������������������       �                     �?�       �                  �&A@+K&:~�?d             c@������������������������       �        ^             b@������������������������       �                     @�       �                   dA�qM�R��?)            �P@������������������������       �                     �?�       �                  �A�U�=���?(            �P@������������������������       �        #            �N@������������������������       �                     @�       K                 �sAg�j�?�          � �@�       D                  ��A�=�0Φ�?�           ��@�       �                   �A��^U���?�           9�@�       �                   ��AП[;U��?&             M@�       �                  R�Ar�qG�?              H@�       �                   *�A�D����?             E@�       �                  ��A�q�q�?             >@�       �                  $\AX�<ݚ�?             2@�       �                  @��@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                  d�A      �?	             (@������������������������       �                     @�       �                  T A      �?              @������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     (@�       �                  D�A�q�q�?	             (@�       �                  @�
AX�<ݚ�?             "@�       �                  h_Aև���X�?             @�       �                   P�A      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   ܗAףp=
�?             $@�       �                  8�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       =                 ,,A&n�VV�?�           �@�                        <�A������?�
           �@�                        DhA�������?�           4�@�                        2A~��t�?�           �@                          �?H>���,�?�           ڧ@������������������������       �        �           �@������������������������       �        �           Đ@                       �:A �>6�t?�            �x@������������������������       �        �            �x@������������������������       �                     �?                        4�Aև���X�?            �A@������������������������       �                     @      	                   �?l��[B��?             =@������������������������       �        
             (@
                       <rA@�0�!��?
             1@������������������������       �                     ,@������������������������       �                     @                       �AL�nIz�?           ��@                       �Ah�˹�?/             S@                       0�A�X�C�?$             L@                         �?H�ՠ&��?#             K@������������������������       �                    �G@������������������������       �                     @������������������������       �                      @������������������������       �                     4@      <                 �GA���0���?�           @�@                        ΥAhǤ���?�           h�@                         �?�(\����?             D@������������������������       �                    �C@������������������������       �                     �?                       DA�j����?�           (�@                       �� A      �?              @������������������������       �                     @                        ��A      �?              @������������������������       �                     �?������������������������       �                     �?       #                 �!�@�96�:�?�           �@!      "                   �?��S�ۿ?             >@������������������������       �                     <@������������������������       �                      @$      1                 �JA������?�           ��@%      *                 �'A(L���?            �E@&      '                 �AX�<ݚ�?             "@������������������������       �                     @(      )                 �8�@z�G�z�?             @������������������������       �                     �?������������������������       �                     @+      .                  ��A�IєX�?             A@,      -                 AA�q�q�?             @������������������������       �                     �?������������������������       �                      @/      0                   �?�g�y��?             ?@������������������������       �                     >@������������������������       �                     �?2      5                 ���@�{��e�?p           ��@3      4                   �?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @6      9                 �eA,��VR��?i           X�@7      8                   �?d��0u��?             >@������������������������       �                     &@������������������������       �        
             3@:      ;                   �?���<��?Y           h�@������������������������       �        �            0x@������������������������       �        ^            @a@������������������������       �        7            �V@>      ?                  ֘A+q�)�?           J�@������������������������       �                     0@@      A                   �?_�w�5�?            :�@������������������������       �        �           b�@B      C                 "IA8�L�$��?c           $�@������������������������       �        �           8�@������������������������       �        t            `g@E      F                   �?N�z���?�            �n@������������������������       �        [             a@G      H                 p�A�C��2(�?D            �[@������������������������       �                    �B@I      J                 �GAd1<+�C�?1            @R@������������������������       �        +            �O@������������������������       �                     $@������������������������       �        a             c@M      t                 lsA���$��?`5          @��@N      O                   �?��*��x?�4          @��@������������������������       �        �           &�@P      a                 ��A R��}F|?.          ��@Q      ^                  ��A pbӪ�>?5*          ���@R      S                  �(A `$���.?*          ���@������������������������       �        �(          @�@T      ]                 0�A�'	�?%           P|@U      \                   �?�a�O�?|            @h@V      W                  D)A g�yB�?Q             `@������������������������       �                     �?X      [                 `��@     ��?P             `@Y      Z                 �l�@@3����?$             K@������������������������       �        #            �J@������������������������       �                     �?������������������������       �        ,            �R@������������������������       �        +            @P@������������������������       �        �            0p@_      `                 lCA �q�q�?             H@������������������������       �                     G@������������������������       �                      @b      c                 ��A���j��?�           `�@������������������������       �                      @d      g                  ��@XLD��?�           X�@e      f                  L�AHm_!'1�??            �X@������������������������       �        :            �V@������������������������       �                      @h      i                  ��A@�S�i��?�           Е@������������������������       �        c           ��@j      o                  |A����O��?-            �Q@k      n                  $�Aףp=
�?             $@l      m                 ��Az�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @p      q                   A����5�?'            �N@������������������������       �                     @r      s                   �?����S��?%             M@������������������������       �                    �D@������������������������       �                     1@u      v                 tiA���x{_�?�            �r@������������������������       �        �            �p@w      �                 ��A     ��?             @@x      y                  ���@l��
I��?             ;@������������������������       �                     @z      �                   �?���|���?             6@{      |                  XA@4և���?             ,@������������������������       �                      @}      �                 ,�Ar�q��?             @~                       �uA      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                 ؍A      �?              @�      �                  F�A      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh~h,h/K ��h1��R�(KM�KK��hJ�Bp      � A    ���@    �R�@     �@    �p�@     ��@     �N@      &@      @      @       @      @       @                      @      �?              M@      @     �A@      @     �@@      @     �@@                      @       @       @       @                       @      7@             R�@     `�@     ��@     `�@     ��@              y@     `�@     �k@      w@             �v@     �k@      @     �k@                      @     `f@     �y@      @              f@     �y@     @W@     �d@     @V@     �d@             �d@     @V@              @             �T@     �n@              7@     �T@     �k@     @R@     `k@             `k@     @R@              $@      @              @      $@             ��@            �D�@     x�@    ��@     �U@    ���@             ؒ@     �U@     Ē@              @     �U@      @      N@             �F@      @      .@       @              @      .@       @       @       @                       @      �?      *@              *@      �?                      ;@    ���@     ��@    ���@     @�@     ��@     @�@     ��@     �{@     ĳ@     @q@     ��@      q@     ��@                      q@      @       @      @                       @     ��@     �d@     ��@                     �d@     ��@     @S@     ��@     �R@              @     ��@      R@     p~@     �C@     p~@                     �C@     �r@     �@@     �r@                     �@@               @     ��@              (@      b@      "@     �V@      @     @T@             @T@      @              @      "@              "@      @              @      K@              K@      @            �A     N�@    H�A    @9�@    РA    ���@     J�@     أ@     s@     �Q@     �h@      F@     �h@      @      ]@      �?      ]@                      �?     @T@      @              �?     @T@      @     @T@                      @              C@      [@      :@     �D@      5@     �D@                      5@     �P@      @     �P@      @      P@       @     �D@              7@       @      *@              $@       @               @      $@              @      �?      @                      �?               @    ���@     L�@     ��@     ��@     ��@     �@     �@      @     �@     �~@     �@                     �~@               @     П@      f@     �u@      3@     �u@                      3@     h�@     �c@     ��@      [@      N@      1@      ?@      ,@      ?@                      ,@      =@      @      =@                      @     ��@     �V@     �J@             ��@     �V@     ��@                     �V@     ��@      I@      f@      @      f@                      @     Px@     �E@               @     Px@     �D@     �v@     �D@     �v@                     �D@      :@                     �U@     ��@     ��@     ��@      j@     ��@                      j@             |�@    �7A    �1�@    � A    �j�@    � A                    �j�@     �@     ȗ@             ��@     �@     �Q@     p{@     �L@     p{@      K@      R@      1@      R@                      1@     �v@     �B@     �s@     �B@     �s@     �A@     �s@     �@@     �q@      9@     �q@                      9@      :@       @      :@                       @       @       @       @                       @               @      J@                      @     �r@      ,@     �m@       @      W@      �?      W@                      �?      b@      @      b@                      @     �N@      @              �?     �N@      @     �N@                      @     ��@     2�@     ��@     ��@     ֦@     �@      :@      @@      1@      ?@      1@      9@      $@      4@      $@       @      �?      @      �?                      @      "@      @      @              @      @      @               @      @              @       @                      (@      @      @      @      @      @      @      �?      @      �?                      @      @                       @      @                      @      "@      �?       @      �?       @                      �?      @             ��@     �@     �@     ֧@     �@     ��@     Ȑ@     ��@     Đ@     �@             �@     Đ@              �?     �x@             �x@      �?              4@      .@      @              ,@      .@              (@      ,@      @      ,@                      @     �g@     ��@      "@     �P@      "@     �G@      @     �G@             �G@      @               @                      4@     �f@     ��@     �f@     �@      �?     �C@             �C@      �?             `f@      }@      @      �?      @              �?      �?              �?      �?             �e@     }@       @      <@              <@       @             @e@     P{@      @     �B@      @      @              @      @      �?              �?      @               @      @@      �?       @      �?                       @      �?      >@              >@      �?             �d@      y@      @       @               @      @             �c@     �x@      3@      &@              &@      3@             @a@     0x@             0x@     @a@                     �V@     8�@     ��@              0@     8�@     ة@             b�@     8�@     `g@     8�@                     `g@      Y@     @b@              a@      Y@      $@     �B@             �O@      $@     �O@                      $@              c@    ���@     �T@    @��@      P@     &�@            ���@      P@    ���@      @     ��@       @    @�@             0|@       @      h@       @     �_@       @              �?     �_@      �?     �J@      �?     �J@                      �?     �R@             @P@             0p@              G@       @      G@                       @     p�@      N@               @     p�@      M@     �V@       @     �V@                       @     �@      I@     ��@              5@      I@      �?      "@      �?      @              @      �?                      @      4@     �D@      @              1@     �D@             �D@      1@             �q@      3@     �p@              *@      3@       @      3@              @       @      ,@      �?      *@               @      �?      @      �?      �?              �?      �?                      @      @      �?      �?      �?      �?                      �?      @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��!XhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B(          f                    �?|ٵ����?;$         ��A       ;                  JHA��z��?��         ��A                          �A�[���P�?(�         HA                          ���@���+���?�f         �^A                           ��@��).�ؓ?�M          ���@                           �?��G����?�M           ��@������������������������       �        &           =�@                           �? ˫�B��?�2          ���@	       
                  xA\k_�l�?!           �@������������������������       �        �            ��@������������������������       �        �            @k@                         :yA�R��Y�?n           l�@������������������������       �        7           �@������������������������       �        7            @U@������������������������       �                     @                           �?@i��J��?8         ��
A������������������������       �        l�          ��@                           �? U�U�ܒ?�]         �GA                          xA@'NH�?��          �r�@������������������������       �        ��          � �@������������������������       �        K           ��@������������������������       �        �z           9�@                           �?� M9Yd�?F!          �{�@                         �xA���A_��?�           ��@������������������������       �        e           N�@������������������������       �        $             N@       8                   ��A���J��?�          �6�@       %                  �+�@P������?           ��@                          �9A��n��?�           ܝ@                           �?�tk~X$�?�           @�@������������������������       �        -           ��@������������������������       �        �           �@!       $                  �7�@�7��?            �C@"       #                    �?�r����?	             .@������������������������       �                     *@������������������������       �                      @������������������������       �                     8@&       -                   �A���}��?I           �@'       *                   ��A�o;����?_            �c@(       )                    �?�sly47�?/            �R@������������������������       �                      J@������������������������       �                     7@+       ,                    �?�L"p�?0            �T@������������������������       �                     B@������������������������       �                    �G@.       /                    �?\�~S/��?�           S�@������������������������       �        Q
           t�@0       3                  ��A@z�J�?�           ��@1       2                  txA ���eK�?{           d�@������������������������       �        j           �@������������������������       �                     4@4       5                  �A���{h�?           `|@������������������������       �                     �?6       7                  �oA �kakd�?           P|@������������������������       �                   `{@������������������������       �                     .@9       :                    �?^F<A�5�?�            Pp@������������������������       �        a            �b@������������������������       �        G            �[@<       M                    �?B���T �?�J          @��@=       >                    �?��aVe��?�           R�@������������������������       �        �           ��@?       L                    �?�:���?           ��@@       G                  ��A�������?           py@A       D                  rA��/�^�?�            �x@B       C                  �mA�C��2(�?             6@������������������������       �                     4@������������������������       �                      @E       F                  �YA0�z��?�?�            @w@������������������������       �        �            �v@������������������������       �                     @H       I                   p�@8�Z$���?
             *@������������������������       �                     @J       K                  �A����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                   x�@N       U                    �?�F,�?B           !�@O       T                    �?࿁�2�?�*          @��@P       S                   n�AԷ�R��?�           ��@Q       R                  BxA�c8�N�?�           \�@������������������������       �        �           �@������������������������       �        8            �U@������������������������       �        �             v@������������������������       �        �          ��@V       e                    �?$���DW�?S          �_�@W       `                  0hA(%�=�P�?J           �@X       [                  �4A�摋���?j             d@Y       Z                   ��A�K�	H�?d             c@������������������������       �        ]            `a@������������������������       �                     ,@\       ]                  �gA      �?              @������������������������       �                     @^       _                  �A���Q��?             @������������������������       �                      @������������������������       �                     @a       d                  �xA�r�6z��?�           Ĩ@b       c                   �A�Lz�<�?�           ~�@������������������������       �        \           8�@������������������������       �        j            `d@������������������������       �                    �A@������������������������       �        	           ��@g       h                    �?�nK�M�u?HQ          ��@������������������������       �        �           �@i       �                   ��A���6���?Z5          @�@j       m                    ��@ p�`�`?3          �-�@k       l                    ��@��"pK�?V            ``@������������������������       �        U            @`@������������������������       �                     �?n       �                    �? 6�K�_?�2           �@o       p                  �zA ���hh?!           .�@������������������������       �        �            ��@q       x                  ܁A8��8���?q             h@r       u                   ���@�X����?             6@s       t                  �qA      �?             (@������������������������       �                     @������������������������       �                     @v       w                  �(Aףp=
�?             $@������������������������       �                     "@������������������������       �                     �?y       |                   P�A`ۘV�?e            @e@z       {                  TA�O4R���?"            �J@������������������������       �        !             J@������������������������       �                     �?}       ~                   WA��-�=��?C            @]@������������������������       �                      @       �                   .A���}<S�?B            �\@�       �                  ��A������?+            �Q@������������������������       �                     4@�       �                  %Aj�q����?             I@������������������������       �                    �D@������������������������       �                     "@�       �                  p�A����?�?            �F@�       �                  �A�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     A@������������������������       �        �           ػ@�       �                  >FA���M@�?M           Ќ@������������������������       �                   p�@�       �                    �?f<t=9%�?B             [@������������������������       �        )            �P@�       �                  ��A�Ń��̧?             E@������������������������       �                    �C@�       �                   �[A�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�bh~h,h/K ��h1��R�(KK�KK��hJ�B0	      �A     ��@    �A     ��@    8A     +�@    (,A     X�@    @<�@      s@    @<�@     �r@     =�@            ���@     �r@     ��@     @k@     ��@                     @k@     �@     @U@     �@                     @U@              @    �d
A     ��@    ��@            �A     ��@    � �@     ��@    � �@                     ��@     9�@             "�@     ն@     N�@      N@     N�@                      N@     ��@     ��@     ̦@     �@     (�@     H�@     �@     ��@             ��@     �@               @     �B@       @      *@              *@       @                      8@     �@     �@     �Q@      V@      7@      J@              J@      7@             �G@      B@              B@     �G@             v�@     ��@             t�@     v�@      B@     �@      4@     �@                      4@     `{@      0@              �?     `{@      .@     `{@                      .@     �[@     �b@             �b@     �[@             ��@    @��@     �x@     8�@             ��@     �x@     Ȋ@     �x@      $@      x@       @      4@       @      4@                       @     �v@      @     �v@                      @      &@       @      @              @       @      @                       @             x�@    ��@    @��@     �@    ���@     �@     `{@     �@     �U@     �@                     �U@              v@            ��@     R�@     ��@     R�@     @k@     �a@      4@     `a@      ,@     `a@                      ,@       @      @              @       @      @       @                      @     8�@     �h@     8�@     `d@     8�@                     `d@             �A@             ��@    ��@      V@     �@            @��@      V@    �(�@      5@     @`@      �?     @`@                      �?     �@      4@     $�@      4@     ��@             �e@      4@      .@      @      @      @      @                      @      "@      �?      "@                      �?     �c@      *@      J@      �?      J@                      �?     @Z@      (@               @     @Z@      $@     �N@      "@      4@             �D@      "@     �D@                      "@      F@      �?      $@      �?      $@                      �?      A@             ػ@             ��@     �P@     p�@             �D@     �P@             �P@     �D@      �?     �C@               @      �?              �?       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJC�NhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaMGhbh,h/K ��h1��R�(KMG��hi�B�G         �                   �AP�C�Â�?y#         ��A       +                  JHA�b��dg�?��         ��A                         �wA@D�q+�?��         t�A������������������������       �        ��         ��A                           �?�S�f�4�?�	           p�@������������������������       �        d           t�@       &                    �?δ� i��?�           ��@       !                   ��@0{�v��?�            pw@	                           �?Hn�.P��?�             o@
                         *�A �#�Ѵ�?i            �e@                         ~�AĴF���?4            �T@                         �}�@ �\���?3            �S@                           �?�θ�?	             *@������������������������       �                     $@������������������������       �                     @                           0�@����e��?*            �P@                         8VA      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        (             P@������������������������       �                     @                           m�@�E�����?5            �V@������������������������       �        /            �S@                         �b�@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@                         ��A�}�+r��?/             S@                           �?`Ql�R�?            �G@������������������������       �                     G@������������������������       �                     �?                            �?ܷ��?��?             =@������������������������       �                     :@������������������������       �                     @"       #                   ��@X�GP>��?R            �_@������������������������       �                      @$       %                    �?ĭ����?Q            @_@������������������������       �        J             \@������������������������       �                     *@'       *                    �?��i���?�           ȡ@(       )                    �?��V�*��?           �@������������������������       �        U           �@������������������������       �        �           (�@������������������������       �        �            �k@,       {                    �?p�ӹ�a�?<O           5�@-       z                    �?`̀��?�           ��@.       Y                  �qA�K�ӫ�?�           l�@/       T                   @y�@��p8�c�?4          ���@0       G                  �}A�q�QQ�?`           ��@1       D                   �@�s��3��?           ��@2       3                  �xAև���X�?            �A@������������������������       �                     @4       A                    Y�@      �?             @@5       <                   `��@�+e�X�?             9@6       7                  �7A�q�q�?	             (@������������������������       �                     @8       ;                   ��@      �?              @9       :                  ���@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @=       @                   ��@8�Z$���?             *@>       ?                   �}@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@B       C                  �YA؇���X�?             @������������������������       �                     @������������������������       �                     �?E       F                    �?$�p���?�           ��@������������������������       �        -           p~@������������������������       �        �            �t@H       I                    �?�N�#/�?Q            @`@������������������������       �        5            �W@J       O                  @�Ab�h�d.�?            �A@K       N                   �~�@X�<ݚ�?             "@L       M                   oAr�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @P       Q                  |A$�q-�?             :@������������������������       �                     ,@R       S                  �cAr�q��?             (@������������������������       �                     $@������������������������       �                      @U       V                    �?@/�̊��?�           b�@������������������������       �                     �?W       X                  �xA`ؠ}o��?�           a�@������������������������       �        �           ��@������������������������       �        C            �X@Z       k                    �?�62���?�           ��@[       f                   ���@��+g��?}             i@\       ]                    �?z�G�z�?y            `h@������������������������       �        \            �b@^       c                   ��@t/*�?            �G@_       `                   �:�@�?�|�?            �B@������������������������       �                     4@a       b                  �AA�IєX�?             1@������������������������       �                     0@������������������������       �                     �?d       e                  �A�z�G��?             $@������������������������       �                     @������������������������       �                     @g       h                  ���@�q�q�?             @������������������������       �                      @i       j                  �XA      �?             @������������������������       �                      @������������������������       �                      @l       w                  $�A����Y�?           `�@m       v                  ��A �w{�t�?           �@n       u                  ��A���ڳ��?j           H�@o       r                    �?@���@�?i           @�@p       q                  �]A ������?�            �w@������������������������       �        �            @w@������������������������       �                     @s       t                   �A��swɃ?            �i@������������������������       �        ~            �i@������������������������       �                     �?������������������������       �                     �?������������������������       �        �             o@x       y                  L�A�c����?           `y@������������������������       �                   �x@������������������������       �                     *@������������������������       �                   ��@|       �                  z�A�(�����?b3           C�@}       �                  (fAXÁu���?V3          �=�@~                           �?��E�B��?7           �@������������������������       �        �           P�@�       �                  `]A@���a��?J            �\@������������������������       �        /            �R@�       �                    �?�(\����?             D@������������������������       �                     "@�       �                  ��A�g�y��?             ?@������������������������       �                     >@������������������������       �                     �?�       �                    B@H���|��?1          @^�@�       �                    �?z�G�z�?             @������������������������       �                      @�       �                    0@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                  ~wA�[[|%��?1           ]�@�       �                    �?h�-%��?m0          @�@�       �                    �?���.��?           �@������������������������       �        [           Ԡ@������������������������       �        �            pp@�       �                    �?���h�h�?j*           ��@������������������������       �        @&          �9�@������������������������       �        *           ��@�       �                  �A�;�=5�?�            0q@�       �                    �?@c��$�?�            �p@������������������������       �                    �D@�       �                   f�A �����?�            @l@�       �                    �?P��`ئ?�            `k@������������������������       �        �            �h@�       �                    �?�GN�z�?             6@������������������������       �                     1@������������������������       �                     @�       �                  �A����X�?             @������������������������       �                      @������������������������       �                     @�       �                  ��A      �?              @������������������������       �                      @������������������������       �                     @�       �                    �?�X����?             6@������������������������       �                     .@������������������������       �                     @�                          �?��n�(��?�(          ��@�       �                    �?vL��4��?�$          ���@�       �                   ��A��>a�?�           г@�       �                  nxA��f��5�?�           ²@�       �                   Z�@X-}�p�?�           x�@�       �                    �?�c�Α�?             =@�       �                   E�@��.k���?             1@�       �                  �xA"pc�
�?
             &@������������������������       �                     "@������������������������       �                      @������������������������       �                     @������������������������       �                     (@�       �                  &�A�ƞ��7�?�           [�@�       �                    �?,�*�?|�?�           <�@�       �                   ��A�t��?P           ��@�       �                  dGA(��4���?O           ��@������������������������       �        �           ��@������������������������       �        �            �n@������������������������       �                      @�       �                  �HA|�n��T�?�           �@������������������������       �        V           ��@������������������������       �        E             Y@�       �                   lVAS*�\�?�           ��@�       �                  xIA,��e�?>           ��@������������������������       �                   Љ@������������������������       �        +            �N@�       �                   pXA �����?q           0�@�       �                   �WA�q�q�?             (@�       �                  �hAև���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?����d��?l           Ё@�       �                  WA��a���?�             w@������������������������       �        �            u@������������������������       �                    �@@�       �                   J�A0w-!��?�             i@�       �                   -A(l58��?            �h@������������������������       �        q            �e@������������������������       �                     9@������������������������       �                     �?������������������������       �        /            �R@�       �                   ��A 7���B�?�            �p@�       �                    �?|�űN�?I            @]@�       �                  H��@�>����?0            @T@�       �                  >GA8�Z$���?             :@������������������������       �                     6@������������������������       �                     @�       �                   �Ah㱪��?!            �K@������������������������       �                     �J@������������������������       �                      @�       �                  ��A�X�<ݺ?             B@������������������������       �                     A@������������������������       �                      @�       �                   ��A`#`��k�?d             c@�       �                  �XA�1���܋?^            @b@������������������������       �        ]             b@������������������������       �                     �?�       �                  dA؇���X�?             @�       �                  @�A�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?�c��o�?           ���@������������������������       �        �           ��@�                        2xAJ(w؏�?�           t�@�       �                   ��A��jL���?g           �@�       �                  GAL�$@t�?�           ��@������������������������       �        D           ؋@������������������������       �        G             _@�       �                   0�@�3���h�?�           &�@�       �                    t@      �?             @������������������������       �                      @������������������������       �                      @�                         0A�.�A�?�           �@�       �                  �fA0�%*�(�?�            pw@�       �                  0��@@3����?c            @d@�       �                  ��@��<D�m�?"            �H@�       �                   lA`Ql�R�?!            �G@������������������������       �                    �D@�       �                   zAr�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �        A            @\@�                        x�Ap���p�?�            �j@�                        ��Aҳ�wY;�?             1@�       �                   2�Ad}h���?
             ,@������������������������       �                     �?                         A8�Z$���?	             *@������������������������       �                     @                        �A�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @                       �0A@9G��?            �h@������������������������       �        {            �g@������������������������       �                      @	      
                 �IA���c&��?�           `�@������������������������       �        |           ��@������������������������       �        q            �e@������������������������       �                     H@                        �A@��NE�?           �@                         �?@�6|���?�             j@                       ��A �w5�?K            �]@������������������������       �        H            �\@                         �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        =            �V@      B                   �? 	|��?           ��@      %                 ��A��&�|�?P           �@                       �gA �	,���?�           x�@                       �KA ��*i?�           P�@������������������������       �        �           (�@                       .[Az�G�z�?             @������������������������       �                     �?������������������������       �                     @      $                 T�A���=�/�?0            @Q@      !                 ��A�n_Y�K�?.            @P@                          �?JJ����?!            �G@������������������������       �                     6@������������������������       �                     9@"      #                   �?r�q��?             2@������������������������       �                     @������������������������       �                     .@������������������������       �                     @&      '                   �?U���y�?�            �m@������������������������       �        2             U@(      )                  x�A؇���X�?Z            @c@������������������������       �                     �?*      -                  �AL紂P�?Y             c@+      ,                 ��A���7�?             F@������������������������       �                     E@������������������������       �                      @.      3                 �#ARԅ5l�??            @[@/      2                  L�Aףp=
�?             $@0      1                  t;Az�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @4      ;                  $zAW�!?�?<            �X@5      8                 pHA�iʫ{�?            �J@6      7                  $5A      �?             @������������������������       �                      @������������������������       �                      @9      :                 :^A؇���X�?            �H@������������������������       �                     E@������������������������       �                     @<      =                  ��A��<b�ƥ?             G@������������������������       �                    �B@>      ?                 �A�����H�?             "@������������������������       �                     @@      A                 ��A�q�q�?             @������������������������       �                      @������������������������       �                     �?C      F                  PA �[oj�?/           �~@D      E                 `0A�����׫?X            �a@������������������������       �        V            `a@������������������������       �                     @������������������������       �        �             v@�t�bh~h,h/K ��h1��R�(KMGKK��hJ�Bp      �A    @��@    |�A    ���@    ��A     |�@    ��A             2�@     |�@     t�@             ��@     |�@      ;@     �u@      (@     �m@       @     �d@      @     �R@      @     �R@      @      $@              $@      @              �?     @P@      �?      �?      �?                      �?              P@      @              �?     @V@             �S@      �?      $@      �?                      $@      @      R@      �?      G@              G@      �?              @      :@              :@      @              .@      \@       @              *@      \@              \@      *@             �@     �@     (�@     �@             �@     (�@             �k@            �0�@    ��@    �+�@     ��@    ���@     ��@     y�@     ��@     �w@     ؂@     �u@     `@      4@      .@              @      4@      (@      3@      @       @      @      @              @      @      @      �?      @                      �?              @      &@       @      �?       @      �?                       @      $@              �?      @              @      �?             �t@     p~@             p~@     �t@              =@     @Y@             �W@      =@      @      @      @      @      �?      @                      �?              @      8@       @      ,@              $@       @      $@                       @     ��@     �X@      �?             ��@     �X@     ��@                     �X@     ��@     `f@     �E@     �c@     �C@     �c@             �b@     �C@       @      B@      �?      4@              0@      �?      0@                      �?      @      @      @                      @      @       @       @               @       @               @       @             �@      5@     Љ@       @     �@       @     �@      @     @w@      @     @w@                      @     �i@      �?     �i@                      �?              �?      o@             �x@      *@     �x@                      *@     ��@             �@    �@�@     �@    �<�@     �\@     X�@             P�@     �\@      �?     �R@             �C@      �?      "@              >@      �?      >@                      �?     D�@     z�@      @      �?       @               @      �?              �?       @             4�@    �y�@     �@    @7�@     pp@     Ԡ@             Ԡ@     pp@             ��@    �9�@            �9�@     ��@              "@     �p@      @     @p@             �D@      @     `k@      @     �j@             �h@      @      1@              1@      @               @      @       @                      @       @      @       @                      @      @      .@              .@      @             ��@     ��@     h�@     W�@     ��@     ��@     ��@     `�@     ��@      ~@      5@       @      "@       @      "@       @      "@                       @              @      (@             ��@     �}@     ��@     �u@     ��@     �n@     ��@     �n@     ��@                     �n@               @     ��@      Y@     ��@                      Y@     ��@      `@     Љ@     �N@     Љ@                     �N@     �@     �P@      @       @      @      @      @                      @              @     �@     �M@     u@     �@@     u@                     �@@     �e@      :@     �e@      9@     �e@                      9@              �?             �R@     @p@      $@     @[@       @     �R@      @      6@      @      6@                      @     �J@       @     �J@                       @      A@       @      A@                       @     �b@       @      b@      �?      b@                      �?      @      �?       @      �?       @                      �?      @             ��@     !�@             ��@     ��@     �v@     ��@     �s@     ؋@      _@     ؋@                      _@     ��@      h@       @       @       @                       @     ��@     �g@     `v@      1@     �c@      @      G@      @      G@      �?     �D@              @      �?              �?      @                       @     @\@             �h@      ,@      &@      @      &@      @              �?      &@       @      @              @       @               @      @                      @     �g@       @     �g@                       @     ��@     �e@     ��@                     �e@              H@     ��@      Q@     �i@      �?     @]@      �?     �\@               @      �?       @                      �?     �V@             ��@     �P@     ��@     �O@     0�@     �D@     H�@      �?     (�@              @      �?              �?      @              =@      D@      9@      D@      6@      9@      6@                      9@      @      .@      @                      .@      @              k@      6@      U@             �`@      6@              �?     �`@      5@      E@       @      E@                       @     �V@      3@      �?      "@      �?      @              @      �?                      @     @V@      $@      F@      "@       @       @       @                       @      E@      @      E@                      @     �F@      �?     �B@               @      �?      @               @      �?       @                      �?     �~@      @     `a@      @     `a@                      @      v@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�R�[hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaMwhbh,h/K ��h1��R�(KMw��hi�BR         &                 xA�-��H5�?"         ��A       {                    �?0>��)��?�         ��A                         NHA�lu�(ܖ?          �`�@������������������������       �        ]�           ��@       V                   �A<��E���?�          ���@       U                    �?�7c���?,           ��@       
                   ܍@��w�{�?�           �@       	                   ���@      �?             (@������������������������       �                     @������������������������       �                     @       P                  B?Ax?��&Y�?�           ��@       O                    �?��X..��?�           ��@       6                    ��@<Sw�[��?�           ��@       -                  @l�@&�w���?)           ~@       ,                   @K�@l������?\            �b@                          ֙@���C�:�?Z            `b@������������������������       �                     �?       '                  �A�M�N���?Y            @b@                         ���@�nkK�?T            @a@                         �N�@�����H�?             ;@                          ���@`2U0*��?             9@������������������������       �        
             4@                         ���@z�G�z�?             @������������������������       �                     @                          ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @       $                  pdA�?�|�?E            �[@                          ���@�L��ȕ?<            @W@������������������������       �        2            @S@        #                  `A      �?
             0@!       "                   �q�@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@%       &                  zoA�����H�?	             2@������������������������       �                      @������������������������       �                     0@(       )                  ��A      �?              @������������������������       �                      @*       +                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @.       3                  �� Aʩ��M��?�            �t@/       2                  p� A�eP*L��?             &@0       1                   ���@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @4       5                    �?�l8ɠ��?�            t@������������������������       �        �            @p@������������������������       �        %            �N@7       L                   ���@PV�,��?�             u@8       K                  |2ADK{22�?�             r@9       H                  TA\2R}�?�            r@:       G                  ��A�F����?b            @c@;       D                  ~2AȨBR��?a             c@<       =                  �� A�X�C�?"             L@������������������������       �                     ?@>       ?                  �A��H�}�?             9@������������������������       �        	             .@@       C                    ��@ףp=
�?             $@A       B                  A      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @E       F                    �? �q�q�??             X@������������������������       �        ;             W@������������������������       �                     @������������������������       �                      @I       J                    �? 7���B�?Q            �`@������������������������       �        M            @`@������������������������       �                     @������������������������       �                     �?M       N                    �?�q�q��?             H@������������������������       �                    �B@������������������������       �                     &@������������������������       �        �           ��@Q       T                    �?�IєX�?�            0t@R       S                    �?��2(&�?             6@������������������������       �                     3@������������������������       �                     @������������������������       �        �            �r@������������������������       �        �	           h�@W       r                  �A@���	H�?w           ��@X       o                   �Ar�q��??            �V@Y       \                  ��A�<p���?:            �T@Z       [                    �?P�Lt�<�?             C@������������������������       �                    �B@������������������������       �                     �?]       l                   V�A"pc�
�?              F@^       i                    �?8����?             7@_       h                   D�A      �?             0@`       g                  �A��
ц��?
             *@a       f                  ƱA�eP*L��?             &@b       c                   ��A����X�?             @������������������������       �                     �?d       e                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @j       k                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?m       n                  ��A���N8�?             5@������������������������       �                     �?������������������������       �                     4@p       q                    �?      �?              @������������������������       �                      @������������������������       �                     @s       v                   ��AzQ����?8           p@t       u                    �?Hm_!'1�?3           �~@������������������������       �                    |@������������������������       �                     D@w       z                  ��
A�n_Y�K�?             *@x       y                    �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @|       �                    �?��,KK��?�         �x	A}       ~                  JHA��v�Wo�?l=           b�@������������������������       �        .7           ��@       �                    �?���z��?>           �@������������������������       �        �           ��@������������������������       �        �             o@�       �                   `�A��8�?%�         �lA�       �                  8HA��_�*�?�         �'A�       �                    �? �u.��
?a         (A�       �                    �? �y���?��          ���@�       �                   �A @�u"?R�          `!�@�       �                   �=A  e��"�>O�          0!�@�       �                   �=A @�s�?H^          @��@������������������������       �        G^           ��@������������������������       �                     �?������������������������       �        �           ��@������������������������       �                     @������������������������       �        {           �@������������������������       �        ��          `��@�       �                  �JA����Ӓ�?�+          @&�@�       �                    �?      �?8             V@�       �                    �?�������?(             N@������������������������       �                      G@������������������������       �                     ,@�       �                    �?����X�?             <@������������������������       �                     4@������������������������       �                      @�       �                    �?��� l�?|+          @�@������������������������       �        '          ���@������������������������       �        `           Л@�       �                  ��A���?           J�@�       �                    �?lJJ�C>�?�           ��@�       �                    �?@��7��?t           ܷ@������������������������       �        �           ��@�       �                  >FA�]l*7��?|           0�@������������������������       �        P           `�@������������������������       �        ,             M@�       �                   "�A��D0�?�           ��@�       �                    �?x2�AGA�?�           H�@�       �                  ��A���8�?           ��@�       �                  8xApbN�;��?!           �@�       �                  �GA� �*+<�?j           ܛ@������������������������       �        �           �@������������������������       �        r            �f@�       �                  *7A���p�?�            �p@������������������������       �        �            p@������������������������       �                     ,@�       �                  0�A�?���?�           ȇ@�       �                  :�A����X�?             @������������������������       �                      @������������������������       �                     @�       �                  pHAlI�
%��?�           ��@�       �                   Z�A|��Y���?�            pu@�       �                  GA�摋���?�             t@������������������������       �        �            �q@������������������������       �                     D@�       �                  NsA�G��l��?             5@������������������������       �                     &@������������������������       �                     $@�       �                  $(Ad��ѩ��?            �y@������������������������       �        �            �w@������������������������       �                    �A@������������������������       �        �            Pr@�       �                   ר@ �=�腱?�            `s@������������������������       �                     �?�       �                    �?��l��?�            Ps@�       �                  �GA/\a��?�            �q@�       �                  
<A�}�+r��?b             c@������������������������       �        Z             b@������������������������       �                      @�       �                   .�A ����?T            @`@�       �                   ��A >��@�?Q            @_@������������������������       �        5            �T@�       �                  HA qP��B�?            �E@�       �                  ��A      �?	             0@������������������������       �                     .@������������������������       �                     �?������������������������       �                     ;@�       �                   \�Az�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     ;@�                        ��A�z�m�,�?           ��@�       �                  ��@R�ѫ��?�           ��@�       �                   ��A؇���X�?             5@�       �                  z�A�}�+r��?             3@������������������������       �                     (@�       �                  ��A؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�                         ��AԄ!K��?�           �@�                          �?f�Sc��?�           p�@�       �                   �#A��,̍S�?�           ��@�       �                  ���@��$
���?�            `s@������������������������       �                      @�       �                  
�AX�Cc�?�            @s@�       �                  4_AX�<ݚ�?i            �f@�       �                    �?~�4_�g�?f             f@������������������������       �        :             Y@������������������������       �        ,             S@������������������������       �                     @�       �                  ��A     ��?Q             `@������������������������       �        
             0@�       �                  .�A���X�?G             \@������������������������       �                     @�       �                    �?���{��?C            @Z@������������������������       �        .            �T@������������������������       �                     7@�       �                   �1A&ᦠ�~�?�            �s@������������������������       �                     <@�       �                  @ �@������?�             r@������������������������       �                      @�                        4�A�E��ӭ�?�             r@�       �                  j�A$Z9��?h            �d@�       �                    �?��h!��?"            �L@������������������������       �                    �D@������������������������       �                     0@�       �                   H>A�2����?F            �[@�       �                  PAA      �?             @�       �                  �`�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                  ��A�����?B            �Z@������������������������       �        	             ,@�       �                  ��AJ� ��w�?9             W@������������������������       �                     �?�                         @�A8�Z$���?8            �V@�       �                   �PA ��~���?7            �V@������������������������       �                     4@�                        ��@z��R[�?,            �Q@                          �?      �?	             $@������������������������       �                     @������������������������       �                     @                       yA�r����?#             N@      	                  �dA�^����?"            �M@                        2\A���|���?             &@������������������������       �                     @                         �?և���X�?             @������������������������       �                     @������������������������       �                     @
                         �?      �?             H@������������������������       �                    �F@������������������������       �                     @������������������������       �                     �?������������������������       �                     �?                         �?|;�p)�?T            @^@������������������������       �        5            �R@������������������������       �                     G@������������������������       �        (             M@                         �?�d�����?             3@                         �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@                       ��A�?�0�!�?S             a@                        ĻA��+7��?	             7@                       �A�KM�]�?             3@                       r�A���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     ,@������������������������       �                     @       !                   �? (��?J            @\@������������������������       �        4            @T@"      %                 "LA     ��?             @@#      $                 6A\-��p�?             =@������������������������       �                     @������������������������       �                     9@������������������������       �                     @'      <                   �?�sr���?u           G�@(      ;                   �? 5�j�?�           �@)      :                 �HA�<��}�?}           l�@*      5                 �Q�@�~_ �?#           $�@+      .                 @��@��D��I�?�            �t@,      -                  �A�nkK�?<             W@������������������������       �        9             V@������������������������       �                     @/      0                 ���@���R��?�             n@������������������������       �        }            �i@1      2                 z�Aг�wY;�?             A@������������������������       �                     9@3      4                   �?�����H�?             "@������������������������       �                      @������������������������       �                     �?6      7                 n�@�'�
��?U           ��@������������������������       �                     @8      9                  4�A,�N��	�?T           ȍ@������������������������       �        0           ȋ@������������������������       �        $             P@������������������������       �        Z            @b@������������������������       �        f            @e@=      d                   �?���}�?�           �@>      ?                   �?p<L�g�?�           Х@������������������������       �        �           ��@@      c                 |�Aƻ�<�5�?D           @�@A      B                   �?��q���?B           0�@������������������������       �        7            �V@C      Z                 f�A���#U��?           X�@D      Y                  ��AH�~�k|�?�           X�@E      V                 n�A��D���?w           �@F      I                  (&�@��Xx��?c           (�@G      H                 .�A�n`���?(             O@������������������������       �        !             I@������������������������       �                     (@J      M                  � A y~.�n�?;           p~@K      L                 �ZAXCږ���?           �z@������������������������       �        
           `y@������������������������       �                     9@N      S                  �*A      �?             L@O      P                  �	A؇���X�?             @������������������������       �                     @Q      R                 h�A�q�q�?             @������������������������       �                      @������������������������       �                     �?T      U                 �|A@�E�x�?            �H@������������������������       �                     H@������������������������       �                     �?W      X                 ��A�q�q�?             >@������������������������       �                     4@������������������������       �                     $@������������������������       �                     D@[      ^                  �AA     p�?}             h@\      ]                 @:A�IєX�?y            `g@������������������������       �        r             f@������������������������       �                     &@_      b                  z�Az�G�z�?             @`      a                 @vA      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @e      l                 �AdP-���?�            �q@f      g                 RMAh��Q(�?)            �P@������������������������       �        !            �I@h      i                 L�A      �?             0@������������������������       �                     &@j      k                  �A���Q��?             @������������������������       �                     @������������������������       �                      @m      t                 �XA �#�Ѵ�?�            �j@n      o                 :�A����?�            �i@������������������������       �        �             i@p      q                  �� Az�G�z�?             @������������������������       �                      @r      s                 A�q�q�?             @������������������������       �                     �?������������������������       �                      @u      v                 ��Aףp=
�?             $@������������������������       �                     "@������������������������       �                     �?�t�b��^     h~h,h/K ��h1��R�(KMwKK��hJ�Bp      D&A    �v�@    �A    �/�@    ��@     ȓ@     ��@            �L�@     ȓ@    �.�@     �@     )�@     �@      @      @              @      @             #�@     ��@     �@      �@     �[@      �@     �S@      y@      (@      a@      $@      a@      �?              "@      a@      @     �`@      @      8@      �?      8@              4@      �?      @              @      �?      �?      �?                      �?       @              @      [@      �?      W@             @S@      �?      .@      �?      @      �?                      @              &@       @      0@       @                      0@      @      @       @              �?      @              @      �?               @             �P@     �p@      @      @      @      @      @                      @      @             �N@     @p@             @p@     �N@              @@      s@      5@     �p@      4@     �p@      .@     `a@      *@     `a@      "@     �G@              ?@      "@      0@              .@      "@      �?      �?      �?      �?                      �?       @              @      W@              W@      @               @              @     @`@             @`@      @              �?              &@     �B@             �B@      &@             ��@              s@      3@      @      3@              3@      @             �r@             h�@              N@     ��@      .@     �R@      "@     @R@      �?     �B@             �B@      �?               @      B@      @      0@      @      $@      @      @      @      @       @      @      �?              �?      @              @      �?              @                       @              @      �?      @              @      �?              �?      4@      �?                      4@      @       @               @      @             �F@     �|@      D@      |@              |@      D@              @       @      @      @              @      @                      @    hzA    @��@    @"�@     ��@     ��@              o@     ��@             ��@      o@             �A    ���@    X;A    ���@    A      @    `��@      @     !�@      @     !�@      �?     ��@      �?     ��@                      �?     ��@                      @     �@            `��@             (�@    ���@      6@     �P@      ,@      G@              G@      ,@               @      4@              4@       @             Л@    ���@            ���@     Л@             ��@     ;�@     ~�@     ��@     `�@     е@             ��@     `�@      M@     `�@                      M@     f�@     pr@     �@     �q@     ƣ@     �q@     �@     @h@     �@     �f@     �@                     �f@     p@      ,@     p@                      ,@     ��@     �V@       @      @       @                      @     �@     @U@     Pr@      I@     �q@      D@     �q@                      D@      &@      $@      &@                      $@     �w@     �A@     �w@                     �A@     Pr@             �r@      &@              �?     �r@      $@      q@      $@      b@       @      b@                       @      `@       @      _@      �?     �T@              E@      �?      .@      �?      .@                      �?      ;@              @      �?              �?      @              ;@             �q@      �@     �p@     �|@      @      2@      �?      2@              (@      �?      @      �?                      @       @             �p@     p{@     �o@      {@     @h@      {@      \@     �h@       @             �[@     �h@      T@      Y@      S@      Y@              Y@      S@              @              >@     �X@              0@      >@     �T@      @              7@     �T@             �T@      7@             �T@     �m@              <@     �T@      j@       @              T@      j@      A@     �`@      0@     �D@             �D@      0@              2@      W@      @      �?      �?      �?      �?                      �?       @              .@     �V@              ,@      .@     @S@      �?              ,@     @S@      *@     @S@              4@      *@     �L@      @      @              @      @               @      J@      @      J@      @      @              @      @      @              @      @              @     �F@             �F@      @              �?              �?              G@     �R@             �R@      G@              M@              ,@      @      �?      @              @      �?              *@              *@     �^@      @      1@       @      1@       @      @              @       @                      ,@      @              @     �Z@             @T@      @      9@      @      9@      @                      9@      @             V�@     8�@     ��@     @k@     �@     @k@     �@      R@     �t@      @      V@      @      V@                      @      n@      �?     �i@             �@@      �?      9@               @      �?       @                      �?     ȋ@     �P@              @     ȋ@      P@     ȋ@                      P@             @b@     @e@              �@     ��@     ��@     T�@             ��@     ��@     @i@     ��@      i@             �V@     ��@     @[@     h�@     �W@     h�@      K@     �@      F@      I@      (@      I@                      (@     p|@      @@     `y@      9@     `y@                      9@     �H@      @      �?      @              @      �?       @               @      �?              H@      �?      H@                      �?      4@      $@      4@                      $@              D@      f@      .@      f@      &@      f@                      &@      �?      @      �?      �?      �?                      �?              @               @      p@      8@     �J@      ,@     �I@               @      ,@              &@       @      @              @       @             �i@      $@     �i@      �?      i@              @      �?       @               @      �?              �?       @              �?      "@              "@      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�v}hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaM�hbh,h/K ��h1��R�(KM���hi�B�_         t                    �?�~�t|�?Y$         ��A       )                  NHA�BS�2�?�         @��@                           �? $��BN?�          `��@������������������������       �        �          ���@                          |�A ����)Q?*�          ���@                          ��@   ?��           ��@                         �A �a/UUE?�           ��@������������������������       �        �           ȧ@	                           �? 7���B�?             ;@
                           �?�}�+r��?             3@                          �KA�X�<ݺ?
             2@������������������������       �        	             1@������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                         �
A �({$M?X�          0<�@                         R�A P�<�%?8w           ��@������������������������       �        �v          ���@                         ��A��V9��?�            �q@������������������������       �                     �?                           �?�#	M���?�            �q@������������������������       �        u            �g@                          ΥAx��B�R�?>            �V@                          ��A }�Я��?<            @V@������������������������       �        :            �T@                          ��Ar�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �         U          `��@       (                    �?�)��OŖ?C	           .�@        #                  H��@���Д^�?X           (�@!       "                  �zA A��� �?i           `�@������������������������       �        d           0�@������������������������       �                     @$       %                   ��A����e��?�           ��@������������������������       �                      @&       '                   wA�{8�?�           ��@������������������������       �        �           H�@������������������������       �                     A@������������������������       �        �            0x@*       K                    �?*���?�           ��@+       .                    �?���
l��?�           ��@,       -                    �?�/ C-��?           ��@������������������������       �        �           X�@������������������������       �        K            �\@/       B                  �wA�	�Q���?�           J�@0       7                   d�@HM����?V           �@1       4                  � A�:�^���?            |@2       3                   uA�LQ�1	�?P            @a@������������������������       �        G             ^@������������������������       �        	             2@5       6                   $�A��)�G��?�            �s@������������������������       �        �             r@������������������������       �                     6@8       =                  ��Axq7.N��?@           (�@9       :                   J�A Q�L�i�?:           �@������������������������       �        f           ζ@;       <                    �?�4�����?�            u@������������������������       �        �            `s@������������������������       �                     ;@>       ?                  �A�<ݚ�?             "@������������������������       �                     �?@       A                   ��A      �?              @������������������������       �                     @������������������������       �                     �?C       F                  z�A@��8��?=             X@D       E                    �?      �?              @������������������������       �                     @������������������������       �                     �?G       H                  ��A�|���?7             V@������������������������       �        0            �S@I       J                    �?ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?L       M                  pHA ��ר�?L
           6�@������������������������       �                      @N       Q                    �?h��|tt�?K
           4�@O       P                  �hA i~z�?0           �~@������������������������       �        ,           ~@������������������������       �                      @R       m                   �A �S��?	           ��@S       b                   �9�@ ��.i\�?�           �@T       a                    �?�1��k�?�             s@U       `                   �-�@�g�y��?�            pq@V       _                  �1A��*����?�            `q@W       Z                   ���@�]��?x            �i@X       Y                  �wA���%yU�?C            �`@������������������������       �        B            ``@������������������������       �                      @[       \                   ���@�F��O�?5            @R@������������������������       �                      @]       ^                  DuA����Q8�?4            �Q@������������������������       �        0            �P@������������������������       �                     @������������������������       �        -             R@������������������������       �                     �?������������������������       �                     9@c       d                  �xA`u�y(�?�           ��@������������������������       �        �           *�@e       j                  ��A�:�]��?            �I@f       i                  >�A��<b�ƥ?             G@g       h                  ��Ar�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     D@k       l                    �?���Q��?             @������������������������       �                      @������������������������       �                     @n       q                  �=A�{�9�?~            `j@o       p                    �?���(\O�?d             d@������������������������       �        Y            �a@������������������������       �                     1@r       s                    �?d,���O�?            �I@������������������������       �                     C@������������������������       �                     *@u       p                 RHA�v�Q���?Z         ��	Av       �                  xAp��6yO�?��         �9Aw       �                    �?��ʻ��?��         �Ax       �                    �?@��ը��?Ǡ         ��Ay       �                  H>A�Eƺ��?�         ��@z       }                    5@X�b)��?d         Ю�@{       |                   �1@�q�q�?             "@������������������������       �                     @������������������������       �                     @~       �                   �`@F݈5��?`         @��@       �                   ``@��G���?            �B@�       �                   �A@؇���X�?            �A@�       �                   �1@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                  h�Aܷ��?��?             =@������������������������       �                     .@�       �                    �?d}h���?             ,@������������������������       �                      @�       �                  ��A      �?             @������������������������       �                      @�       �                   �_@      �?             @�       �                  �wA      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                  ~A`p����?G         ��@�       �                  �A�@�C�гʸ?�          ��@�       �                    �?�a=�1n�?�6          @��@������������������������       �        }           Z�@�       �                  ��@�6)r��?~0           +�@�       �                   P�A�v��u^�?10          ��@������������������������       �        ]-          ���@������������������������       �        �           ��@�       �                  �"�@�Y>J��?M            @]@�       �                  $�A��.k���?
             1@������������������������       �                     @�       �                   �@A"pc�
�?             &@������������������������       �                      @������������������������       �                     "@�       �                   r�A0w-!��?C             Y@������������������������       �        9            �U@������������������������       �        
             *@�       �                   �A�Ll�Z�?�          �Q�@������������������������       �        ��           M�@������������������������       �        n
           G�@�       �                  JAx�iЬ�?J	           ��@�       �                  iAP`���?	           
�@�       �                    �?l����?�           0�@������������������������       �        �            �s@�       �                   ؐA ��b��?$           ��@������������������������       �        �           <�@������������������������       �        ~            �g@�       �                   ؖA�y5�w�?%           h�@������������������������       �                   X�@������������������������       �                     A@�       �                  j/Ar�q��?-             R@�       �                  )Aև���X�?	             5@�       �                   ��Ar�q��?             (@������������������������       �                     $@������������������������       �                      @�       �                   A�<ݚ�?             "@������������������������       �                      @������������������������       �                     @�       �                    �?�IєX�?$            �I@������������������������       �                     $@�       �                  |AA��p\�?            �D@�       �                  .�A"pc�
�?             &@������������������������       �                     @�       �                  �@A�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                  �A(;L]n�?             >@�       �                  t�A      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     <@�       �                   "�A�摋���?f             d@������������������������       �        ]            �a@������������������������       �        	             4@������������������������       �        ��           ��@������������������������       �        �.          ���@�       �                   ،@w�e��?           f�@������������������������       �                     @�       �                  f~A�������?           X�@�       �                   �s�@����_�?y             h@�       �                  pA�C��2(�?             6@������������������������       �                     3@�       �                  `~A�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   ƌA�\��N��?l            `e@�       �                    �?"�!���?i            �d@�       �                   ��A:%�[��?Y            �a@�       �                   �.�@8^s]e�?9            �U@�       �                    �?      �?             >@������������������������       �        
             .@������������������������       �                     .@�       �                  z|A���y4F�?'            �L@�       �                  �{A�d�����?             C@�       �                    �?r�q��?             >@������������������������       �                     9@������������������������       �                     @�       �                  2|A      �?              @�       �                  |A      �?             @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                   P	A�KM�]�?             3@������������������������       �                      @�       �                    �?"pc�
�?             &@������������������������       �                     "@������������������������       �                      @�       �                  �yA\�����?             �K@������������������������       �                     @�       �                    �?���H.�?             I@������������������������       �                     5@������������������������       �                     =@������������������������       �                     9@������������������������       �                     @�       O                   �?�,^�~o�?�           ֤@�                         ��@�jq3��?Q           l�@�       �                   ���@ I��� �?�           ��@������������������������       �        "             O@�       �                    �?��8����?_           ��@�       �                    �?|E+�	��?o            @d@������������������������       �        f            �b@������������������������       �        	             *@�                        l�A`�zE�0�?�            Pw@�       �                   �P�@@�0�!��?             A@�       �                   P�@r�q��?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�                         Z�Ah�����?             <@������������������������       �                     4@                       ��A      �?              @������������������������       �                     �?������������������������       �                     @                       ���@ (��?�            0u@                       ���@�H�I���?H            @\@������������������������       �        9            �U@      
                 ��A ��WV�?             :@      	                  �5�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     7@                         �?�=|+g��?�            @l@������������������������       �        �            �i@������������������������       �                     4@      D                 \/AåI$`�?�           �@      ;                 �
A�VRA<�?�           ��@                        (��@�T�����?�           h�@������������������������       �                      @      "                 45A�F��I�?�           X�@                        (R A��e���?i           h�@                        d% A      �?             @������������������������       �                      @                        �G A      �?             @                       ̼A      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                       ���@��	�
�?d           8�@                         �?�(�ڡ)�?�            0w@������������������������       �        �            �s@������������������������       �        $            �K@       !                   �? �h�7W�?|            �j@������������������������       �        s             i@������������������������       �        	             (@#      (                 dA��[�p�?7            �W@$      '                 QA"pc�
�?             &@%      &                   �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @)      6                 D�A�o��gn�?3            �T@*      /                  L�A¦	^_�?             ?@+      .                  ��A�C��2(�?
             &@,      -                  ,�Az�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @0      1                  �GA���Q��?	             4@������������������������       �                     @2      3                  ��A�t����?             1@������������������������       �                     @4      5                 0�A�q�q�?             (@������������������������       �                     @������������������������       �                     @7      :                  ��A ��WV�?              J@8      9                   �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                    �G@<      ?                  	AX�<ݚ�?             2@=      >                  hXAz�G�z�?             $@������������������������       �                      @������������������������       �                      @@      C                  ʦA      �?              @A      B                   �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?E      L                 �AI��M��?#           p|@F      I                 �A�a�� �?�             m@G      H                   �?85�}C�?J            �^@������������������������       �        C             \@������������������������       �                     $@J      K                   �?Ц�f*�?F            �[@������������������������       �        C            �Z@������������������������       �                     @M      N                   �?X�*��?�            �k@������������������������       �        �            `h@������������������������       �                     <@P      k                 ��AF�k��V�?C           ��@Q      j                 �A�e鷎r�?"           ��@R      W                  p��@�_��y�?           x�@S      V                 ��A�DÓ ��?F            @Y@T      U                   �?<���D�?E            �X@������������������������       �        >            �U@������������������������       �                     (@������������������������       �                      @X      i                   �?H��ԛ�?�           P�@Y      f                 ��A���7�?�           ��@Z      ]                 f�AX����4�?�           P�@[      \                  �A���IBk�?�           `�@������������������������       �        ~           Ȃ@������������������������       �                     3@^      a                 �Ar�q��?             >@_      `                  �\Az�G�z�?             @������������������������       �                     �?������������������������       �                     @b      e                 4A`2U0*��?             9@c      d                  �A      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     5@g      h                 6�A���Q��?             $@������������������������       �                     @������������������������       �                     @������������������������       �        %             K@������������������������       �                    �@@l      o                  PA     ��?!             P@m      n                  4�@8�Z$���?             J@������������������������       �                      @������������������������       �                     F@������������������������       �                     (@q      r                   �?h'¡��?�5           A�@������������������������       �        0          ��@s      �                 *sA��yDv�?�           l�@t      u                   �?м{��$�?i            �@������������������������       �        �            �q@v      �                 ��A�K(v��?�           ȝ@w      �                   �?�Abe�?�           d�@x      �                 4�A ܼ!f�?a           �@y      �                 ��A���C��?>            �Z@z      {                 ���@,���j�?=            �Y@������������������������       �                     >@|      �                 6oA0�й���?,            @R@}      �                 �A@�E�x�?            �H@~                       �3A �q�q�?             8@������������������������       �                     7@������������������������       �                     �?������������������������       �                     9@�      �                  ��A�q�q�?             8@������������������������       �                     0@������������������������       �                      @������������������������       �                     @�      �                 F�A���U�?#           ��@�      �                 �A�H�G�հ?!           ��@������������������������       �        ?             X@�      �                  �APu�?�           ��@������������������������       �        �           ��@������������������������       �                     =@�      �                  �PA�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        V           ��@�      �                   �?��9��Ϸ?           �y@�      �                 �A4��6�?�            Pp@�      �                 �+A@�0�!��?*             Q@�      �                 (?A`�Q��?             9@�      �                 �zA��s����?             5@������������������������       �                     @�      �                 ��A������?	             .@������������������������       �                      @�      �                  �YA8�Z$���?             *@������������������������       �                     &@������������������������       �                      @������������������������       �                     @�      �                 tA�ʈD��?            �E@�      �                  znAև���X�?             @������������������������       �                     @������������������������       �                     @�      �                 d�A������?             B@������������������������       �                    �@@�      �                 @	A�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                  ��A(�f+�W�?|             h@������������������������       �        w             g@������������������������       �                      @������������������������       �        ]            �b@�      �                 ��A>A�F<�?             C@�      �                  
A4?,R��?             B@�      �                   �?HP�s��?             9@������������������������       �                     7@������������������������       �                      @�      �                  4�A���!pc�?             &@�      �                  �dA      �?             @�      �                 `�A      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�t�bh~h,h/K ��h1��R�(KM�KK��hJ�BP      �A    ���@    PX�@     ��@    p��@     �G@    ���@            ���@     �G@    ���@      @     ��@      �?     ȧ@              :@      �?      2@      �?      1@      �?      1@                      �?      �?               @            �;�@      @    ���@      @    ���@             `q@      @              �?     `q@      @     �g@              V@      @      V@      �?     �T@              @      �?              �?      @                       @    `��@             ڬ@      E@     ԩ@      E@     0�@      @     0�@                      @     H�@      B@               @     H�@      A@     H�@                      A@     0x@             �@      �@     ��@     $�@     �\@     X�@             X�@     �\@             ��@     �{@     ��@      v@     �y@      D@      ^@      2@      ^@                      2@      r@      6@      r@                      6@     �@     �s@     �@     `s@     ζ@              ;@     `s@             `s@      ;@              @       @              �?      @      �?      @                      �?       @     �W@      �?      @              @      �?              �?     �U@             �S@      �?      "@              "@      �?             ~�@     �n@               @     ~�@     �n@     ~@       @     ~@                       @     ��@     �m@     ��@      L@     pr@      "@     �p@      "@     �p@       @     �h@       @     ``@       @     ``@                       @     �P@      @               @     �P@      @     �P@                      @      R@                      �?      9@             2�@     �G@     *�@              @     �G@      �?     �F@      �?      @      �?                      @              D@      @       @               @      @              >@     �f@      1@     �a@             �a@      1@              *@      C@              C@      *@             �A     v�@    8PA     -�@    �/A     �@    8�A     �@    �W�@     �@    O�@     ��@      @      @      @                      @    �N�@     ��@      >@      @      >@      @      @       @      @                       @      :@      @      .@              &@      @       @              @      @               @      @      �?      �?      �?              �?      �?               @                       @    �L�@     �@    �n�@     �@    ���@     ��@     Z�@            ���@     ��@    ���@     ��@    ���@                     ��@     �W@      6@       @      "@      @               @      "@       @                      "@     �U@      *@     �U@                      *@     M�@     G�@     M�@                     G�@     ��@     �m@     H�@      l@     ��@     �g@     �s@             <�@     �g@     <�@                     �g@     X�@      A@     X�@                      A@      N@      (@      (@      "@      $@       @      $@                       @       @      @       @                      @      H@      @      $@              C@      @      "@       @      @              @       @      @                       @      =@      �?      �?      �?      �?                      �?      <@             �a@      4@     �a@                      4@     ��@            ���@             X�@     t�@      @             <�@     t�@     �T@     �[@       @      4@              3@       @      �?              �?       @             @T@     �V@     @T@     �U@      L@     �U@      ;@      N@      .@      .@              .@      .@              (@     �F@      $@      <@      @      9@              9@      @              @      @      @      @      @      �?              �?      @                       @       @               @      1@               @       @      "@              "@       @              =@      :@              @      =@      5@              5@      =@              9@                      @     ��@     ��@     �f@     ��@      D@     h�@              O@      D@     �~@      *@     �b@             �b@      *@              ;@     �u@      @      <@      @      �?      @               @      �?              �?       @              �?      ;@              4@      �?      @      �?                      @      5@     �s@      �?      \@             �U@      �?      9@      �?       @               @      �?                      7@      4@     �i@             �i@      4@             �a@     ȏ@      Y@     ؂@      W@     ��@       @             �V@     ��@     �Q@     8�@      @      @               @      @      �?      �?      �?              �?      �?               @             �P@      �@     �K@     �s@             �s@     �K@              (@      i@              i@      (@              4@     �R@      "@       @      @       @               @      @              @              &@      R@      "@      6@      �?      $@      �?      @              @      �?                      @       @      (@      @              @      (@              @      @      @              @      @               @      I@       @      @              @       @                     �G@       @      $@       @       @       @                       @      @       @      @      �?              �?      @                      �?     �D@     �y@      *@     `k@      $@      \@              \@      $@              @     �Z@             �Z@      @              <@     `h@             `h@      <@             8�@      a@     ؆@     @]@     Ѕ@     @]@      ,@     �U@      (@     �U@             �U@      (@               @             `�@      >@     ��@      >@     ��@      8@     Ȃ@      3@     Ȃ@                      3@      9@      @      �?      @      �?                      @      8@      �?      @      �?      @                      �?      5@              @      @      @                      @      K@             �@@              F@      4@      F@       @               @      F@                      (@     ��@    �*�@            ��@     ��@     @W@     ��@      O@     �q@             М@      O@     ��@      E@     ��@      E@     �W@      (@     �W@      "@      >@              P@      "@      H@      �?      7@      �?      7@                      �?      9@              0@       @      0@                       @              @     ȉ@      >@     ��@      =@      X@             ��@      =@     ��@                      =@       @      �?       @                      �?     ��@             Px@      4@      n@      4@      L@      (@      1@       @      1@      @      @              &@      @               @      &@       @      &@                       @              @     �C@      @      @      @      @                      @     �A@      �?     �@@               @      �?       @                      �?      g@       @      g@                       @     �b@              @      ?@      @      ?@       @      7@              7@       @              @       @      @      �?      �?      �?      �?                      �?       @                      @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg}�XhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaMShbh,h/K ��h1��R�(KMS��hi�B(J                           :�A\؋^%v�?�#         ��A                          ���@�S�j�?:�         ��A                         pHA���5A��?_          @��@                           �? F(b5��?pU          ���@������������������������       �        �          ���@                          ��@ �QQ���?�7          ��@                         xA���0SI�?�7          ��@������������������������       �        �6          @��@	       
                    �?��0�?�            �u@������������������������       �        �            �s@������������������������       �                     <@                          ��@      �?             @������������������������       �                     @������������������������       �                     �?                           �?�/[y�e�?�	           ڮ@                         8_A�"�V�J�?C           �@                           �?��n2An�?4           ��@                           �?��H�}�?�           \�@������������������������       �        �           ��@������������������������       �                   pz@������������������������       �        _             c@������������������������       �                     8@                           �?��ϷJ�?k           L�@������������������������       �        �           :�@                           ��@ �����?�            �p@                         ��AP���Q�?             4@������������������������       �                     3@������������������������       �                     �?                         �jA���n��?�            �n@������������������������       �        �            �n@������������������������       �                     �?        �                    �?@�D����?�         ��A!       H                    �?L�8t�m�?�W         ��A"       #                  {A �t��Qj?R�          ���@������������������������       �        r�          @Y�@$       9                   r�@�d�n8�?�           X�@%       ,                  r�AH.�!���?>             Y@&       )                  p�A��S���?
             .@'       (                  �A����X�?             @������������������������       �                     @������������������������       �                      @*       +                  XKA      �?              @������������������������       �                      @������������������������       �                     @-       8                   k�@P�;�&��?4            @U@.       5                    �?���O1��?3            �T@/       2                  j�Ar�q��?             K@0       1                   ���@ 7���B�?             ;@������������������������       �                     �?������������������������       �                     :@3       4                  d�Al��
I��?             ;@������������������������       �        	             3@������������������������       �                      @6       7                  �Aܷ��?��?             =@������������������������       �                     :@������������������������       �                     @������������������������       �                      @:       ?                    �?���I�?�           Ȑ@;       <                  ({A���ym�?�            �@������������������������       �                      @=       >                  �HA�ޛ(���?�           �@������������������������       �        �           �@������������������������       �        *            @P@@       C                   <�A��h��?�            �t@A       B                  48A��\m���?�            �i@������������������������       �        r             e@������������������������       �                    �B@D       E                   6MA@���|N�?Y             `@������������������������       �                    �A@F       G                  �]A�*/�8V�?D            �W@������������������������       �        <             U@������������������������       �                     $@I       V                   z�Aج�<o�?E�         HQAJ       M                  �wAOX��?[`         �cAK       L                  HHA�Ֆ���?[         @ A������������������������       �        +7         ���@������������������������       �        �#          �w�@N       U                  Z0A&�Ǹ���?U           �@O       R                  ��A�{�}:�?�           ��@P       Q                    �?�C�ݳ"�?�           О@������������������������       �        8           �@������������������������       �        �           ��@S       T                    �?�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �        q            �f@W       �                  �{Ady�l��?�&          ���@X       �                   r�A�U�w/��?V&           a�@Y       �                  ���@��8"��?�           ��@Z       }                  @�@��
�8B�?!           0~@[       b                   �A,���j�?�            �i@\       ]                   ڋA���N8�?             5@������������������������       �        
             *@^       _                   :�A      �?              @������������������������       �                     @`       a                   ��A���Q��?             @������������������������       �                     @������������������������       �                      @c       |                  ���@�f����?z             g@d       {                   ��A���.�6�?y             g@e       v                  ��@�˹�m��?d             c@f       i                    �?,�T�6�?F             Z@g       h                  `�At�e�í�?*            �P@������������������������       �        '             O@������������������������       �                     @j       o                   ��@�MI8d�?            �B@k       l                   x�@ 7���B�?             ;@������������������������       �                     3@m       n                  \�A      �?              @������������������������       �                     @������������������������       �                     �?p       q                   ��A      �?	             $@������������������������       �                      @r       s                   �A      �?              @������������������������       �                     @t       u                   ~�A      �?             @������������������������       �                     @������������������������       �                     �?w       z                    �?@��8��?             H@x       y                  ��A�?�|�?            �B@������������������������       �                     B@������������������������       �                     �?������������������������       �                     &@������������������������       �                     @@������������������������       �                     �?~                         ��A�?}<�%�?�            Pq@������������������������       �        �            q@������������������������       �                     @�       �                    �?�ۊ��+�?�           6�@�       �                  :HA���yR�?           ̜@������������������������       �                   (�@������������������������       �        i             e@�       �                  �SA4�[���?3           @�@������������������������       �        �           Ј@������������������������       �        4            �S@�       �                   ��A��^�@G�?�           "�@������������������������       �                     @�       �                   �|@�DT��;�?�          � �@�       �                   �t@�eP*L��?             &@�       �                   �Z@r�q��?             @�       �                   ��A      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �w@z�G�z�?             @������������������������       �                      @�       �                  �!A�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?��$Y+�?y           �@�       �                   VA�8���
�?�           ]�@�       �                  ���@(L���?�           ��@������������������������       �                     E@�       �                  V0A��e�1�?�           0�@������������������������       �        ^           0�@������������������������       �        3             X@�       �                   d%Al��G�?#           ��@�       �                  �#A�==Q�P�?�            �q@������������������������       �        �            @q@������������������������       �        	             "@�       �                  ���@k���?}           ��@�       �                  nGA^��8�?�           2�@������������������������       �        )           ��@������������������������       �        �            �h@�       �                   �%A$w7��+�?�           w�@�       �                  lA�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   �@H�+>�?�           q�@�       �                   ��A      �?             (@�       �                   dAև���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   ��A𭐇���?�           e�@�       �                  �JAl���k#�?o           �@������������������������       �        D
           �@������������������������       �        +           �|@�       �                   ��AD����\�?X            ``@������������������������       �                     @�       �                  �-A�J�4�?V            @_@�       �                  p�A��s����?J            @Z@�       �                   |�Ar�q��?H            �Y@�       �                   ԏAr٣����?1            �P@�       �                  hoAf1r��g�?(            �J@�       �                   D�A �o_��?             9@�       �                  �1A؇���X�?             ,@������������������������       �                     (@������������������������       �                      @�       �                  #A�eP*L��?	             &@������������������������       �                     @�       �                   �A      �?              @������������������������       �                     @�       �                  huA      �?             @������������������������       �                     @������������������������       �                     �?�       �                  ��Ah�����?             <@������������������������       �                     ;@������������������������       �                     �?�       �                   8�A�n_Y�K�?	             *@������������������������       �                     @�       �                   �AX�<ݚ�?             "@������������������������       �                     @�       �                  ��A�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   ��A������?             B@������������������������       �                    �A@������������������������       �                     �?������������������������       �                     @������������������������       �                     4@�       �                   Z�A�QEܡg�?�
           ٰ@�       �                   B�A��Q �?�
           ��@�       �                   d�APa�	�?C            �X@�       �                  vHA�KM�]�?             3@������������������������       �                     1@������������������������       �                      @�       �                   h�A@�z�G�?1             T@������������������������       �        %             P@�       �                  jqA      �?             0@������������������������       �                     .@������������������������       �                     �?�       �                   b�A�q�Bw�?J
           M�@������������������������       �                     @�       �                  "OAlZ��U�?I
           J�@������������������������       �        A	           F�@������������������������       �                   pz@�       �                  �&A���?            �D@������������������������       �                     ?@������������������������       �                     $@�       �                   A|��Q_�?�            `m@�       �                    �?����?|            �i@������������������������       �        L            �\@������������������������       �        0            �V@������������������������       �                     >@�       �                   �rA ��b.�W?�D           �@�       �                   HrA ����b?�           ��@�       �                  �\A ��?_?�           ��@������������������������       �                   Z�@�       �                  d^A���L!��?�           �@������������������������       �                      @�       �                  �pA�����2�?�           �@�       �                  ��A�˹�m��?             C@������������������������       �                    �A@������������������������       �                     @�       �                    �?��W��D�?�           p�@�       �                  �yA� ta��?�           Ȇ@������������������������       �        �           ��@�       �                  Z�Ar�q��?             @�       �                   ��A�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �        �            0x@������������������������       �                      @                        ��A �M�vN?�*          ���@������������������������       �        #*          @��@                       (�Aj���?m             e@������������������������       �                     �?                       �IA �q�q�?l             e@                       ��A�=
ףp�?f             d@������������������������       �        I            �\@      
                  $�A��<b�ƥ?             G@      	                  �A���N8�?             5@������������������������       �                     4@������������������������       �                     �?������������������������       �                     9@                       ��A      �?              @������������������������       �                     @������������������������       �                      @      8                 �HAfh­N��?�(          ���@                         �?���^FU�?�$          ���@                         �?�XNr��?�          ���@                         �?@�{*��?�           H�@                       nxA��b�h�?�           ��@������������������������       �        �           J�@������������������������       �                    �D@������������������������       �        �            `u@                       �:A�>~%���?^           �@                         �?2b��?R           ߷@������������������������       �        �           ��@������������������������       �        s           ؁@                         �?�q�q�?             2@������������������������       �                     (@������������������������       �                     @      #                  ��A�����a�?�           �@      "                  p�A���!5��?m            `f@       !                 �hA@]����?l            @f@������������������������       �        i            �e@������������������������       �                     @������������������������       �                     �?$      7                   �? 1l�£�?@           U�@%      2                 ��A�6�ɹu�?           ��@&      )                   �?��K���?�           �@'      (                 �}A@sV yɉ?S           ��@������������������������       �        M           h�@������������������������       �                     @*      +                  ��A �4����?�           <�@������������������������       �        �            �q@,      /                 �D�@ f}�'6�?�           Ș@-      .                 f~A�Qv���x?�           ��@������������������������       �        �           ��@������������������������       �                      @0      1                 �tA�T�~`��?W            �@������������������������       �        P           ��@������������������������       �                     "@3      4                  N�A     ��?            �@������������������������       �        �            �p@5      6                 �zA �y�ƺ�?l           ̕@������������������������       �        \           d�@������������������������       �                     :@������������������������       �        ,           0}@9      L                   �?Hu�|�?           X�@:      ;                 �k�@� �Q�f�?�           �@������������������������       �        D            �W@<      =                 ��@�[��m&�?b            �@������������������������       �                     @>      ?                   �?ȥ6�?�?a           ��@������������������������       �        %            �@@      E                 �cA���Q��?<            �W@A      D                 �vA��Hg���?            �F@B      C                   �?��>4և�?             <@������������������������       �                     &@������������������������       �                     1@������������������������       �                     1@F      K                  ��Az�):���?              I@G      J                  r�A�[�IJ�?            �G@H      I                   �?      �?             D@������������������������       �                     4@������������������������       �                     4@������������������������       �                     @������������������������       �                     @M      N                   �?P��L��?n           ��@������������������������       �        H           ��@O      R                  �A ������?&            �O@P      Q                 �aA$�q-�?             *@������������������������       �                     (@������������������������       �                     �?������������������������       �                     I@�t�bh~h,h/K ��h1��R�(KMSKK��hJ�B0      , A    @��@    <�A    ���@    `2�@     Ϊ@    ���@      t@    ���@            ���@      t@    @��@     �s@    @��@              <@     �s@             �s@      <@              �?      @              @      �?             0�@     N�@     ��@     @�@     ��@     ��@     pz@     ��@             ��@     pz@              c@                      8@     pp@     >�@             :�@     pp@       @      3@      �?      3@                      �?     �n@      �?     �n@                      �?    ��A    �p�@     uA    �k�@     ��@      a@    @Y�@             8�@      a@     �S@      6@      @       @      @       @      @                       @       @      @       @                      @     �Q@      ,@     �Q@      (@     �F@      "@      :@      �?              �?      :@              3@       @      3@                       @      :@      @      :@                      @               @      �@     �\@     �@     �P@               @     �@     @P@     �@                     @P@     �q@     �G@      e@     �B@      e@                     �B@     �]@      $@     �A@              U@      $@      U@                      $@    (A    �I�@    @��@     T�@    ���@    �w�@    ���@                    �w�@     ؅@     �@     ؅@     �@     ��@     �@             �@     ��@               @      �?              �?       @                     �f@     ��@     ��@    �i�@     ��@     �@     �p@     �|@      6@     �g@      2@      0@      @      *@              @      @              @      @       @      @                       @     �e@      *@     �e@      (@     �a@      (@     @W@      &@      O@      @      O@                      @      ?@      @      :@      �?      3@              @      �?      @                      �?      @      @       @              @      @              @      @      �?      @                      �?     �G@      �?      B@      �?      B@                      �?      &@              @@                      �?     q@      @     q@                      @     H�@     �n@     (�@      e@     (�@                      e@     Ј@     �S@     Ј@                     �S@     ��@     ��@              @     ��@     |�@      @      @      @      �?      �?      �?      �?                      �?      @              �?      @               @      �?       @      �?                       @     ��@     h�@     :�@     �@     ��@      X@      E@             0�@      X@     0�@                      X@     �@     �@     @q@      "@     @q@                      "@     ָ@     Ѕ@     ��@     �h@     ��@                     �h@     ��@     0@       @      @       @                      @     ��@     �~@      @      "@      @      @              @      @                      @     �@     `~@     �@     �|@     �@                     �|@     @Z@      :@              @     @Z@      4@     @U@      4@     @U@      1@      I@      0@     �F@       @      2@      @      (@       @      (@                       @      @      @      @              @      @              @      @      �?      @                      �?      ;@      �?      ;@                      �?      @       @              @      @      @      @               @      @       @                      @     �A@      �?     �A@                      �?              @      4@             D�@     p{@     �@     �z@      X@      @      1@       @      1@                       @     �S@      �?      P@              .@      �?      .@                      �?     F�@     �z@              @     F�@     pz@     F�@                     pz@      ?@      $@      ?@                      $@     �V@      b@     �V@     �\@             �\@     �V@                      >@     �@      4@     ��@      (@     ��@      $@     Z�@             �@      $@               @     �@       @     �A@      @     �A@                      @     \�@      @     ��@      @     ��@              �?      @      �?       @               @      �?                      @     0x@                       @    ���@       @    @��@              d@       @              �?      d@      @     �c@      �?     �\@             �F@      �?      4@      �?      4@                      �?      9@               @      @              @       @             ��@     7�@    ���@     
�@     x�@     ٵ@     ��@     �D@     J�@     �D@     J�@                     �D@     `u@             �@     ��@     ؁@     ��@             ��@     ؁@              @      (@              (@      @             ׳@     �H@     �e@      @     �e@      @     �e@                      @              �?     *�@     �E@     W�@     �E@     �@      1@     h�@      @     h�@                      @     �@      &@     �q@             ��@      &@     ��@       @     ��@                       @     ��@      "@     ��@                      "@     ��@      :@     �p@             d�@      :@     d�@                      :@     0}@             @Z@     ��@     �E@     \�@             �W@     �E@     ȍ@      @              C@     ȍ@              �@      C@     �L@      &@      A@      &@      1@      &@                      1@              1@      ;@      7@      ;@      4@      4@      4@      4@                      4@      @                      @      O@     ��@             ��@      O@      �?      (@      �?      (@                      �?      I@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ	�tlhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaM�hbh,h/K ��h1��R�(KM���hi�B�i         �                    �?�X�3fX�?�#         ��A       M                    �? B1@c�?{         ���@                           �?@�P�]�?]�          @�@                         �HA�YI���?�          ��@������������������������       �        �           �@                           �? ����?           (�@������������������������       �        �           H�@������������������������       �        @             W@	       ,                   ��A �jlm�?��          ���@
                         N�A e �x�e?��          ���@                          @��@ ����"?�          �F�@                         ��A Z���_?�           ,�@������������������������       �        �           �@                          � �@r�q��?             @������������������������       �                     @������������������������       �                     �?                         J�A �
�̯?_�          @��@������������������������       �        Z�          ���@                          P6A�䞠�l�?           �|@������������������������       �        �            �w@                         ��A@�)�n�?-            @U@������������������������       �                     @������������������������       �        ,            �T@                         p�A@�0k�q�?�           Z�@������������������������       �                     �?                         BxA��%���?�           Y�@                          n�A ��<hY8?u           �@������������������������       �        t           �@������������������������       �                     �?                          H0A�5U��K�?8            �T@������������������������       �                    �C@        %                  ��A"pc�
�?             F@!       "                   >A      �?             @@������������������������       �                     3@#       $                   TA$�q-�?             *@������������������������       �                     �?������������������������       �                     (@&       )                  ��A�q�q�?             (@'       (                   ��A؇���X�?             @������������������������       �                     @������������������������       �                     �?*       +                  �Az�G�z�?             @������������������������       �                     �?������������������������       �                     @-       :                  �xA̹�"���?-	           |�@.       /                   �A�-�&b��?
	           �@������������������������       �                      @0       5                   ��A� ����?		           �@1       4                    �?H������?�           v�@2       3                  BAl%<���?�           �@������������������������       �                    ��@������������������������       �        �            �r@������������������������       �        �            ps@6       9                    �?���yv��?o           0�@7       8                  �>A��n/:ֽ?G           �@������������������������       �        4           0~@������������������������       �                     @@������������������������       �        (            �P@;       B                  8lA0B��D�?#            �M@<       ?                  �R�@�S����?             C@=       >                    �?����X�?	             ,@������������������������       �                     $@������������������������       �                     @@       A                    �?�8��8��?             8@������������������������       �                     6@������������������������       �                      @C       L                  LMAև���X�?             5@D       K                  �A�	j*D�?             *@E       F                  ��AX�<ݚ�?             "@������������������������       �                     @G       H                   �A�q�q�?             @������������������������       �                      @I       J                  ��A      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @N       e                  �GA�g�1(Y�?b           u�@O       `                   �A 4��K?�W          @o�@P       Q                  �~A �nƛ2D?�W           l�@������������������������       �        �V          `7�@R       [                  i�@ ���?           `z@S       T                  lA,(��?M            �_@������������������������       �                     �?U       Z                    �? ,V�ނ�?L            �_@V       W                  �A���"�?F             ]@������������������������       �                     7@X       Y                   �yA rpa�?5            @W@������������������������       �        2             V@������������������������       �                     @������������������������       �                     $@\       ]                   ��AP����?�            pr@������������������������       �        �            r@^       _                  ��Ar�q��?             @������������������������       �                     @������������������������       �                     �?a       b                  ��A�J�4�?             9@������������������������       �                      @c       d                   ��A���}<S�?             7@������������������������       �                     5@������������������������       �                      @f       g                  pHA��؂F�??
           .�@������������������������       �                     @h       k                    �?��ٝ���?=
           +�@i       j                  �zA �5yy�?7            @������������������������       �        3           �~@������������������������       �                     @l       �                   �A����Uƾ?	           v�@m       �                    �?@�l�_�?|           Ϊ@n       �                  R�A ;��⧜?�           8�@o       t                  �LA`�~qՙ?X           <�@p       s                   ���@�����?             5@q       r                  �JA�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     2@u       |                  ,GA ;�̫��?K           �@v       y                   H>�@ *;L]n�?�           ��@w       x                  ,vA��k����?�             j@������������������������       �        �             i@������������������������       �                     @z       {                  ZyA`1	��ә?m            �@������������������������       �        [           �@������������������������       �                     <@}       ~                   8tA /���m?V           H�@������������������������       �        �            `v@       �                   6~A@�����?~            `h@������������������������       �                     �?������������������������       �        }            @h@�       �                  ��A���N8�?L            �_@������������������������       �                     �?�       �                  �A`2U0*��?K            @_@������������������������       �        H             ^@������������������������       �                     @������������������������       �        �            �t@�       �                  J�A����&��?�            �j@�       �                    �?Ĝ�oV4�?u            �f@������������������������       �        i             d@������������������������       �                     6@������������������������       �                     >@�       �                  �Ax�E�]�?          �	A�       �                  �wA�< �9�?��         ��A�       �                    �?�}��P�?H�         �*A�       �                    �?�o� j`�?�=         �e�@�       �                  <HAlc s���?�         p+�@������������������������       �        ��          PH�@������������������������       �                   �@������������������������       �        !           ��@�       �                    �?w�Y4�?N�          @��@�       �                  �&�@$3�$�T�?ݙ          �p�@�       �                  �-�@4z�HJp�?�           ��@�       �                  |HA���\��?�           ��@������������������������       �        �           ��@������������������������       �        ?            �X@�       �                    �d@����M��?�           ��@������������������������       �                     @�       �                  KA�U��t�?�           ��@������������������������       �        M           }�@������������������������       �        W           ��@�       �                   ~�A��(Н��?D�          `�@�       �                   `;�@���ӈ�?4�           �@�       �                   �7�@U7��=�?4           "�@�       �                  .�@�U�O���?2           �@�       �                  p��@(�s���?a             e@�       �                  �	�@��pBI�?,            @R@�       �                  rnA���}<S�?             7@������������������������       �                     5@������������������������       �                      @������������������������       �                     I@�       �                  �FA<����?5            �W@������������������������       �        0            �U@������������������������       �                      @�       �                  JJA ;�F��?�           ʢ@������������������������       �                   v�@������������������������       �        �            �r@������������������������       �                     @�       �                   �YAD�w�rY�? �          ���@�       �                  �GA�g��m�?��           ��@������������������������       �        ut          ���@������������������������       �        *           ٴ@�       �                   bA(N"�߾?a           ��@������������������������       �        5             S@�       �                  �]A�J哿�?,           0}@������������������������       �                    {@������������������������       �                    �A@�       �                  �2�@��}*_��?             ;@������������������������       �                      @�       �                   T�A�\��N��?             3@�       �                   �A"pc�
�?             &@�       �                  8+A      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                  �RA      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �        q           �@�       �                   @��@�[V[0�?h           ��@�       �                  ��A)G�� �?           �z@�       �                  D�A��B�5��?�            0p@�       �                  &�A4�^o�]�?K            @\@�       �                    �?f1r��g�?F            �Z@�       �                    �?��<b�ƥ?=             W@������������������������       �        &            �L@�       �                   0��@ >�֕�?            �A@������������������������       �                    �@@������������������������       �                      @������������������������       �        	             ,@�       �                    �?����X�?             @�       �                  �[�@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?���;QU�?a            @b@�       �                    �? 
�V�?X            �`@������������������������       �        >             W@�       �                    �?�Ń��̧?             E@������������������������       �                    �D@������������������������       �                     �?�       �                  ҒA      �?	             (@�       �                  �Aև���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                  ��A�IєX�?b            @e@�       �                    �? �й���?+            @R@������������������������       �        *             R@������������������������       �                     �?�       �                    �?�$��y��?7            @X@������������������������       �        1             V@������������������������       �                     "@�       {                 �FAd[�z�z�?Z           ��@�       (                 B�A½xaSI�?�           ��@�       '                   �?J�����?�           ��@�       �                  `l�@v���?�           ��@�       �                  �M�@�������?             A@������������������������       �                     $@�       �                  @�@      �?             8@�       �                    �@��.k���?             1@������������������������       �                      @�       �                   �A��S���?             .@�       �                   �g�@����X�?             @������������������������       �                      @������������������������       �                     @�       �                  @1�@      �?              @������������������������       �                     @�       �                  �A���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�                         �@Ѓs˛�?�           ��@�                        ��A������?;            �Y@�                        P_AR�����?/             T@�                         yAh�����?             L@�                           �?D�n�3�?             C@������������������������       �                     6@������������������������       �        
             0@                       ��Ar�q��?             2@                         �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     $@      
                 �<A      �?             8@      	                   �?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?                       Z�A�n_Y�K�?             *@                       ��Az�G�z�?             @������������������������       �                     @������������������������       �                     �?                         �?      �?              @������������������������       �                     @������������������������       �                     �?                         �?�LQ�1	�?             7@������������������������       �                     @������������������������       �        	             4@                        �lA��SZ��?\           P�@                       (A�k],=~�?           �{@                         �?��R��?           `{@������������������������       �        �            pp@������������������������       �        i            �e@������������������������       �                     "@      "                 n�A�8~��?A            �Z@                       @��@�uw\l��?8            @W@������������������������       �        
             *@                       ��@      �?.             T@������������������������       �                     @       !                   �?���y4F�?-             S@������������������������       �        "             N@������������������������       �                     0@#      &                 ��Aև���X�?	             ,@$      %                 ��Az�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �        :            �X@)      *                  �6�@DW�T��?�           �@������������������������       �                     @+      0                 �@�@By��ǅ�?�           ̘@,      /                   �?ү�~�?W           ��@-      .                   �?$���?�             v@������������������������       �        �             s@������������������������       �                     I@������������������������       �        w            @g@1      N                 �	A8��
��?�           \�@2      E                  ���@��
n��?�            �q@3      4                 ��A��.k���?             �I@������������������������       �                      @5      8                  � �@�lg����?            �E@6      7                   �?      �?              @������������������������       �                     @������������������������       �                     @9      D                  ��@">�֕�?            �A@:      C                   �?�t����?             A@;      B                 J�Aд>��C�?             =@<      A                  `��@؇���X�?             <@=      >                   T�@����X�?             ,@������������������������       �                     "@?      @                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             ,@������������������������       �                     �?������������������������       �                     @������������������������       �                     �?F      M                   �?���Q��?�            `m@G      J                 ��Ah�����?�             l@H      I                   �?      �?             4@������������������������       �                     $@������������������������       �                     $@K      L                   �?f�B���?            �i@������������������������       �        `            `d@������������������������       �                    �D@������������������������       �                     &@O      n                  ��An �b��?�           ȇ@P      m                   �?��r��,�?�           ��@Q      j                  8A4��.�<�?           p}@R      e                 ��A<\����?           �{@S      V                 ЧA������?�            w@T      U                   �?X'"7��?B             [@������������������������       �        ?            �Y@������������������������       �                     @W      ^                 ��AȰi�o��?�            Pp@X      [                  �
A���|���?             6@Y      Z                 ʰA�8��8��?	             (@������������������������       �                     &@������������������������       �                     �?\      ]                   �?�z�G��?             $@������������������������       �                     @������������������������       �                     @_      b                 .�A=�J�C�?�            �m@`      a                   �?�|����?�            `m@������������������������       �        �            �j@������������������������       �                     5@c      d                   �?      �?             @������������������������       �                      @������������������������       �                      @f      g                  eA��
���?+            �R@������������������������       �                     G@h      i                   �? 	��p�?             =@������������������������       �                     ;@������������������������       �                      @k      l                   �?�+$�jP�?             ;@������������������������       �                     6@������������������������       �                     @������������������������       �        �            �k@o      v                 L�A�xGZ���?-            �Q@p      u                   �?V������?            �B@q      t                 H�A8�Z$���?
             *@r      s                   �?      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     8@w      z                   �?���|���?            �@@x      y                   �?���7�?             6@������������������������       �                     5@������������������������       �                     �?������������������������       �        
             &@|      }                   �?<��ٵ�?�            �o@������������������������       �        �            `j@~      �                  �dA�D����?             E@      �                 ��AP����?             C@�      �                  |cA     ��?             @@�      �                   �?ҳ�wY;�?	             1@������������������������       �                     &@������������������������       �                     @�      �                 0~A��S�ۿ?	             .@������������������������       �                     �?������������������������       �                     ,@������������������������       �                     @������������������������       �                     @�      �                   �?VǤ����?j          ���@�      �                 b,A�I�H��?�          �
�@�      �                  ��A�UcA�,�?k           �@�      �                   �?P�%f��?�           ��@������������������������       �                   Y�@�      �                 @>A@!��{�?�           ��@�      �                  �gA`�I����?|           С@�      �                 @"A� W�{�?�           Н@�      �                  ��@���$/�?u           x�@�      �                 �.Aг�wY;�?&             Q@������������������������       �        %            �P@������������������������       �                      @�      �                 ЈA���ٙ��?O           Ў@������������������������       �        L           ��@������������������������       �                     @�      �                  �A�ܱ�|F�?           ��@�      �                 VdA�_�wd�?R           Ȁ@������������������������       �        J           @�@������������������������       �                     1@�      �                 ��A@ux�ᭉ?�            �s@������������������������       �        �            �s@������������������������       �                      @�      �                 �zA�F�sɪ?�            @w@������������������������       �        �            �v@������������������������       �                     $@�      �                 jAT(y2��?G            �]@������������������������       �        B            �[@������������������������       �                      @�      �                 �hA�T�j��?�           ��@�      �                  ʣ@d�`��8�?�           <�@�      �                  b�A8�Z$���?             *@�      �                  ��A���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�      �                   �?�uw�?�           �@������������������������       �        �           �@������������������������       �        �            �@������������������������       �                     ;@�      �                  ~�A�J'��)�?           ��@�      �                  0�AX;��?7            @V@������������������������       �        6            �U@������������������������       �                     @�      �                  ҘA@Vהf��?H           Ќ@�      �                 X�A ܖ�DRv?�           ��@�      �                 <�A�Ր�m�?           �x@�      �                  ��@��r���t?           �x@�      �                   �? J���#�?�             f@������������������������       �        W            �]@�      �                 @��@0�)AU��?*            �L@������������������������       �        )             L@������������������������       �                     �?������������������������       �        �            �k@������������������������       �                     �?������������������������       �        �            �t@�      �                  ��A�eGk�T�?o            �g@������������������������       �                     �?�      �                  ��@��S����?n            �g@�      �                  �A qP��B�?            �E@�      �                 ���@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                    �@@������������������������       �        T            @b@�      �                 LA�:FձW�?�           ��@�      �                 �^�@������?u           �@�      �                  ��A��s����?             5@�      �                 �qA����X�?	             ,@������������������������       �                     $@������������������������       �                     @������������������������       �                     @�      �                  "A�������?e           p�@�      �                 reA�s��;�?�            @v@������������������������       �        �            Pu@�      �                 4
A���Q��?             .@�      �                  �A"pc�
�?	             &@������������������������       �                     �?�      �                 �Aףp=
�?             $@�      �                 L~A      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                 fIA��C�)&�?�           P�@������������������������       �        V           8�@�      �                   �?��y�:�?*            �P@������������������������       �                    �F@������������������������       �                     6@�      �                 l�A������?             1@������������������������       �                     *@������������������������       �                     @�t�b�W�      h~h,h/K ��h1��R�(KM�KK��hJ�B0      �"A    ���@    �g�@     Ȗ@    @��@     ��@     N�@     H�@     �@              W@     H�@             H�@      W@            ���@     p|@    ���@     @T@     F�@      @     (�@      �?     �@              @      �?      @                      �?    ���@      @    ���@             �|@      @     �w@             �T@      @              @     �T@             �@     @S@              �?     �@      S@     �@      �?     �@                      �?       @     �R@             �C@       @      B@      �?      ?@              3@      �?      (@      �?                      (@      @      @      @      �?      @                      �?      �?      @      �?                      @     ��@     `w@     r�@     �t@               @     r�@     �t@     &�@     �r@     ��@     �r@     ��@                     �r@     ps@             0�@      @@     0~@      @@     0~@                      @@     �P@              .@      F@      @      @@      @      $@              $@      @               @      6@              6@       @              "@      (@      "@      @      @      @      @               @      @               @       @       @               @       @              @                       @    �T�@      p@    `m�@      .@    �j�@      &@    `7�@             �y@      &@     @^@      @              �?     @^@      @     �[@      @      7@              V@      @      V@                      @      $@              r@      @     r@              �?      @              @      �?              5@      @               @      5@       @      5@                       @     v�@     `n@              @     v�@      n@     �~@      @     �~@                      @     ��@     @m@     v�@      F@     �@      F@     �@      C@      3@       @      �?       @      �?                       @      2@             ʦ@      B@     z�@     �A@      i@      @      i@                      @     �@      <@     �@                      <@     @�@      �?     `v@             @h@      �?              �?     @h@              ^@      @              �?      ^@      @      ^@                      @     �t@              6@     �g@      6@      d@              d@      6@                      >@     �A     ?�@    @A    ���@    ��A    @��@    p��@     �@    PH�@     �@    PH�@                     �@     ��@             ��@     ��@    @Z�@     ��@     -�@     ��@     ��@     �X@     ��@                     �X@     }�@     ��@              @     }�@     ��@     }�@                     ��@    �T�@     >�@    �R�@     4�@     ��@     �s@     ��@     @s@     �c@      $@     �Q@       @      5@       @      5@                       @      I@             �U@       @     �U@                       @     v�@     �r@     v�@                     �r@              @    `7�@     ��@    ���@     ٴ@    ���@                     ٴ@     �@     �A@      S@              {@     �A@      {@                     �A@      1@      $@       @              "@      $@       @      "@       @       @       @                       @              @      @      �?              �?      @             �@             ��@     (�@     �D@     @x@      ?@     �l@      5@      W@      0@     �V@       @     �V@             �L@       @     �@@             �@@       @              ,@              @       @      �?       @      �?                       @      @              $@      a@      �?     �`@              W@      �?     �D@             �D@      �?              "@      @      @      @      @                      @      @              $@      d@      �?      R@              R@      �?              "@      V@              V@      "@             �@     �@     ��@     h�@      x@     `y@     �q@     `y@      9@      "@      $@              .@      "@       @      "@               @       @      @       @      @       @                      @      @       @      @              @       @               @      @              @             @p@     �x@     �L@      G@     �B@     �E@      ?@      9@      0@      6@              6@      0@              .@      @      @      @              @      @              $@              @      2@      �?      $@              $@      �?              @       @      @      �?      @                      �?      �?      @              @      �?              4@      @              @      4@             `i@     �u@     �e@      q@     �e@     pp@             pp@     �e@                      "@      <@     �S@      4@     @R@              *@      4@      N@      @              0@      N@              N@      0@               @      @       @       @       @                       @              @     �X@             ��@      �@      @             x�@      �@     �m@      s@      I@      s@              s@      I@             @g@             0x@     ��@     �U@      i@      8@      ;@       @              0@      ;@      @      @              @      @              &@      8@      $@      8@      @      8@      @      8@      @      $@              "@      @      �?              �?      @                      ,@      �?              @              �?              O@     �e@     �I@     �e@      $@      $@              $@      $@             �D@     `d@             `d@     �D@              &@             �r@     �|@     pp@     �z@     �E@     �z@      C@     `y@      B@     �t@      @     �Y@             �Y@      @              ?@     �l@       @      ,@      �?      &@              &@      �?              @      @              @      @              7@      k@      5@     �j@             �j@      5@               @       @               @       @               @     @R@              G@       @      ;@              ;@       @              @      6@              6@      @             �k@              C@      @@      :@      &@       @      &@       @      @              @       @                      @      8@              (@      5@      �?      5@              5@      �?              &@              1@     �m@             `j@      1@      9@      *@      9@      @      9@      @      &@              &@      @              �?      ,@      �?                      ,@      @              @             8�@     M�@     �@     �@     ��@     #�@     h�@     ��@             Y�@     h�@     �E@     ��@     �A@     l�@      9@     `�@      @     �P@       @     �P@                       @     ��@      @     ��@                      @     �@      3@     @�@      1@     @�@                      1@     �s@       @     �s@                       @     �v@      $@     �v@                      $@     �[@       @     �[@                       @     X�@     |�@     X�@     �@      &@       @      @       @      @                       @       @              �@     �@             �@      �@                      ;@      @     `�@      @     �U@             �U@      @              @     ��@       @     І@       @     �x@      �?     �x@      �?     �e@             �]@      �?      L@              L@      �?                     �k@      �?                     �t@       @     �g@      �?              �?     �g@      �?      E@      �?      "@              "@      �?                     �@@             @b@     ��@      O@     H�@      M@      1@      @      $@      @      $@                      @      @             ��@      K@     �u@      "@     Pu@              @      "@       @      "@      �?              �?      "@      �?      �?      �?                      �?               @      @             �@     �F@     8�@              6@     �F@             �F@      6@              *@      @      *@                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ޡhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaM_hbh,h/K ��h1��R�(KM_��hi�B�L                          BHApˎ��`�?�#         ��A       9                  BxA .�6/8�?��         ��A       8                    �? �)�с�?M�         P�A       	                   �A@��u��?�}         h�A                         xA  1�L�>�\          �A������������������������       �        �\         ��A                           �?      �?              @������������������������       �                     @������������������������       �                      @
       /                  ��AB��Xq/�?�           ���@                          õ@��C% �?�           G�@                           �?����O��?~            �j@������������������������       �        0            �T@                           �?��؇>��?N            @`@������������������������       �        -            �O@������������������������       �        !            �P@       .                    �?j}�z)�?          ���@                          B�Adcá�K�?�           ��@                           �?Z�Oy�+�?.           6�@������������������������       �        �           :�@������������������������       �        f           ��@       +                   B�A�-����?�             i@                          R�A�Q����?h             d@������������������������       �                     @       (                  ��@�����?f            �c@                         (��@`��}3��?!            �J@                           �?      �?              @������������������������       �                     �?������������������������       �                     @                          Z�A�<ݚ�?            �F@������������������������       �                     �?        %                   (�@�������?             F@!       $                  �A      �?             0@"       #                    �?�eP*L��?             &@������������������������       �                     @������������������������       �                     @������������������������       �                     @&       '                    �? �Cc}�?             <@������������������������       �                     9@������������������������       �                     @)       *                    �?.y0��k�?E             Z@������������������������       �                    �F@������������������������       �        (            �M@,       -                    �?�G�z�?             D@������������������������       �                     *@������������������������       �                     ;@������������������������       �        n
           ��@0       7                    �? LTC��?1           ��@1       4                  H�A�9�����?o           Ё@2       3                    �?���df�?%           �|@������������������������       �        U            @_@������������������������       �        �            �t@5       6                    �?      �?J             \@������������������������       �                     E@������������������������       �        /            �Q@������������������������       �        �            Pr@������������������������       �        �H          ���@:       �                    �?:|�B1�?e
           ��@;       B                    �?҉����?�           
�@<       A                    �?ȕ�ޡK�?N           ��@=       >                    �?/Ru���?           ��@������������������������       �        8            @W@?       @                   �A��8{�~�?�           ��@������������������������       �        �           h�@������������������������       �                     C@������������������������       �        A            �Y@C       �                  ��Ap�xP{�?e           ��@D       K                    �?<	O�X��?*           (�@E       H                  ��A�s�c���?�            �l@F       G                    �?z�G�z�?3            �V@������������������������       �        *             R@������������������������       �        	             2@I       J                    �?`�q�0ܴ?Y            �a@������������������������       �        U            �`@������������������������       �                     @L       Y                  �AP8Ձ��?�           ��@M       T                  ��A/rX���?           �y@N       O                   P�@h�{�\��?           py@������������������������       �                      @P       S                  �A�$�����?           Py@Q       R                    �?\s�n��?
           0y@������������������������       �        �            0v@������������������������       �        "             H@������������������������       �                      @U       V                  �Aև���X�?             @������������������������       �                     @W       X                    �?      �?             @������������������������       �                     @������������������������       �                     �?Z       �                  $�A`�o�|��?�           �@[       �                  ZA�mؐ���?            ��@\       c                   �2A��R}�v�?�           ��@]       `                   ��@�UM���?�            �w@^       _                   ��@      �?              @������������������������       �                     �?������������������������       �                     �?a       b                    �?�3�ނ��?�            �w@������������������������       �        �            �v@������������������������       �        
             (@d       i                   �At��%�?�            �u@e       f                  �a�@d}h���?"             L@������������������������       �                     �?g       h                    �?z�G�z�?!            �K@������������������������       �                     F@������������������������       �                     &@j                         X��@��� @�?�            r@k       t                  2�A ���g=�?)            @Q@l       m                  ��A��+7��?             7@������������������������       �                     &@n       s                  ��@      �?             (@o       p                   N_A      �?              @������������������������       �                     @q       r                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @u       z                   �A�nkK�?             G@v       y                  `��@r�q��?             @w       x                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @{       ~                  �g�@�(\����?             D@|       }                    �?��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?������������������������       �                     9@�       �                  H�A�2�~w�?�            �k@�       �                  4�A��hJ,�?             A@�       �                    �?@4և���?             <@������������������������       �                     :@������������������������       �                      @�       �                  �A      �?             @������������������������       �                      @�       �                   ��A      �?             @������������������������       �                     �?������������������������       �                     @�       �                  \�AH��2�?y            @g@�       �                    �?`Y����?Z             a@������������������������       �        W            �`@������������������������       �                     @�       �                  ��A i���t�?            �H@������������������������       �                      @�       �                   J�A=QcG��?            �G@�       �                  ��A�Ń��̧?             E@������������������������       �                     C@�       �                  xKA      �?             @������������������������       �                     �?������������������������       �                     @�       �                  �A���Q��?             @�       �                  ��A�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                  �At/*�?9            �W@�       �                  ��A      �?
             0@�       �                   ȹA���!pc�?             &@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                  ��A��-�=��?/            �S@�       �                   �@
AZՏ�m|�?            �H@�       �                   8�@P���Q�?             4@�       �                  ҙAr�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             ,@�       �                  �A>���Rp�?             =@������������������������       �                     "@�       �                  ��A��Q��?             4@������������������������       �                     $@�       �                  ȣA�z�G��?             $@������������������������       �                     @�       �                  RA      �?             @�       �                   ��A      �?             @������������������������       �                      @�       �                  D�A      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     =@�       �                    �?x��r��?�            `j@������������������������       �        z            `g@������������������������       �                     8@�       �                    �?�+e�X�?;             Y@������������������������       �        /             S@������������������������       �                     8@�       �                    �?`�דD�?�           P�@�       �                  B�A��N*tt�?4           `@�       �                  �~A $i���?%           �}@�       �                   @�A�����H�?             B@������������������������       �                     @@������������������������       �                     @�       �                  �A@H�>���?           �{@�       �                    �?x�}���?�            �t@�       �                  �A��"�O��?�            �r@�       �                  N�A8q���?�            �r@�       �                   *�A ���|�?�            Pr@������������������������       �        �            �q@������������������������       �                     "@�       �                   JqA����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     =@������������������������       �        D             [@�       �                   L�A8�Z$���?             :@������������������������       �                     6@������������������������       �                     @�       �                    �?h&��)�?~           x�@�       �                    �@�KM�]�?B            �\@�       �                  ¥A4և����?A             \@�       �                    M�@Hn�.P��?"             O@�       �                  <�A�q�q�?             @�       �                  �A�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                  �:A�h����?             L@������������������������       �                    �H@�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                  ��A�:pΈ��?             I@�       �                  N�A�q�q�?
             .@�       �                  ��Ar�q��?             (@������������������������       �                     �?�       �                  R�A�C��2(�?             &@������������������������       �                     @�       �                  �Az�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                  ��A >�֕�?            �A@�       �                    �?      �?             @@������������������������       �                     ?@������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�                         �A`1��[�?<           `�@�       �                   _AhX�ptE�?           ؊@�       �                   @�Al��?I           ��@������������������������       �        >           p�@�       �                  J�A@4և���?             ,@������������������������       �        	             (@�       �                  ܵA      �?              @������������������������       �                     �?������������������������       �                     �?�       �                  pA0`%w�?�            �s@������������������������       �                      @�                          �?�a-SF�?�            �s@                         ��AL��n��?�            Pr@������������������������       �        �            �p@������������������������       �                     :@������������������������       �                     8@������������������������       �        -            @T@      6                   �?8���g��?�R          �g�@      %                  �A��~���?)           �@                         �?���c�?�          ���@                       BxA��r
'��?�           V�@	                         �?���l��?�           �@
                         �?#_2�?�           Ј@������������������������       �        �            �@������������������������       �        F            �]@������������������������       �        �           Ѹ@                         �? 5x ��??            �Z@������������������������       �        =             Z@������������������������       �                     @                       ��A e'�qƖ?�	           B�@                       ~A�d���?�	            �@������������������������       �        s	           ��@                       ��AP���Q�?             D@                         �? ���J��?            �C@������������������������       �                     C@������������������������       �                     �?������������������������       �                     �?                         J�@�nkK�?\             d@                        p�@�q�q�?             (@������������������������       �                     @������������������������       �                     @                         fqA@m����?W            �b@                       lyA 
�V�?P            �`@������������������������       �        O            �`@������������������������       �                     �?!      $                   �?��S�ۿ?             .@"      #                 �A$�q-�?             *@������������������������       �                     (@������������������������       �                     �?������������������������       �                      @&      3                  ��A`�H�/��?_           ��@'      ,                  NA��:����?[           @�@(      )                  !Aև���X�?             @������������������������       �                      @*      +                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @-      0                 v At���Ú�?X           �@.      /                   �?p�/E�f�?y            �g@������������������������       �        j            �d@������������������������       �                     5@1      2                   �?���偛�?�            Pv@������������������������       �        �            �t@������������������������       �                     6@4      5                   �?�����H�?             "@������������������������       �                     �?������������������������       �                      @7      J                   �?�>���V�?�5          �E�@8      ;                  @m@ CT��c�?W           �@9      :                   �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?<      =                   �?T��?T           �@������������������������       �        �           ��@>      C                   ��@�!��b�?�            0p@?      @                   �?�}�+r��?             3@������������������������       �                     @A      B                 IA$�q-�?             *@������������������������       �                     (@������������������������       �                     �?D      I                  ���@@v�����?�             n@E      H                   �?�Ru߬Α?K            �\@F      G                 �\A�e���@�?3            @S@������������������������       �        2             S@������������������������       �                     �?������������������������       �                    �B@������������������������       �        S            �_@K      R                  ��Apm2�?i/          @��@L      M                   �?��;�	�?�,           ��@������������������������       �        1(           ��@N      O                 {A�.g�4;�?�           x�@������������������������       �                   �@P      Q                   �?|��?���?             ;@������������������������       �                     ,@������������������������       �                     *@S      T                   �?|��ا�?�           ��@������������������������       �        g           �@U      V                 �uA҆�s��??             Z@������������������������       �                      @W      X                   �?r�q��?<             X@������������������������       �        %            �L@Y      Z                 A��-�=��?            �C@������������������������       �                     9@[      ^                  �MA����X�?             ,@\      ]                 ��Aև���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�t�bh~h,h/K ��h1��R�(KM_KK��hJ�B�      ,"A    @��@    x]A     ϼ@     7A     Ե@    ��A     Ե@    ��A       @    ��A              @       @      @                       @     �@     ҵ@     O�@     ?�@     �b@     �O@     �T@             �P@     �O@             �O@     �P@             ��@      �@     ��@      �@     :�@     ��@     :�@                     ��@     @X@     �Y@      U@      S@      @             @T@      S@      B@      1@      �?      @      �?                      @     �A@      $@              �?     �A@      "@      $@      @      @      @      @                      @      @              9@      @      9@                      @     �F@     �M@     �F@                     �M@      *@      ;@      *@                      ;@     ��@             �|@     0y@     �d@     0y@     @_@     �t@     @_@                     �t@      E@     �Q@      E@                     �Q@     Pr@            ���@             <�@     �@     ��@     X�@     ��@      C@     P�@      C@     @W@             h�@      C@     h�@                      C@     �Y@             �g@     ��@     �d@     ��@      8@     �i@      2@      R@              R@      2@              @     �`@             �`@      @             �a@     T�@      L@     `v@      J@     0v@       @              I@     0v@      H@     0v@             0v@      H@               @              @      @      @              �?      @              @      �?             �U@     x�@      O@     ��@      G@     0�@      *@     �v@      �?      �?              �?      �?              (@     �v@             �v@      (@             �@@     �s@      (@      F@      �?              &@      F@              F@      &@              5@     �p@       @     �N@      @      1@              &@      @      @       @      @              @       @      �?              �?       @              @               @      F@      �?      @      �?       @               @      �?                      @      �?     �C@      �?      ,@              ,@      �?                      9@      *@     �i@      @      =@       @      :@              :@       @              @      @       @              �?      @      �?                      @       @     @f@      @     �`@             �`@      @              @      F@       @              @      F@      �?     �D@              C@      �?      @      �?                      @       @      @       @      �?              �?       @                       @      0@     �S@       @       @       @      @      @      @              @      @              @                      @       @     �Q@       @     �D@      �?      3@      �?      @      �?                      @              ,@      @      6@              "@      @      *@              $@      @      @      @              @      @      @      �?       @              �?      �?      �?                      �?               @              =@      8@     `g@             `g@      8@              8@      S@              S@      8@             ��@     �d@      ~@      6@     �|@      2@      @@      @      @@                      @     �z@      ,@     �s@      ,@     r@      ,@     r@      &@     �q@      "@     �q@                      "@      @       @      @                       @              @      =@              [@              6@      @      6@                      @     x�@     �a@      (@     �Y@      $@     �Y@      @     �M@       @      @       @      �?       @                      �?              @      �?     �K@             �H@      �?      @              @      �?              @     �E@      @      $@       @      $@      �?              �?      $@              @      �?      @      �?                      @      @               @     �@@      �?      ?@              ?@      �?              �?       @               @      �?               @             �@     �D@     ��@     �D@     x�@      *@     p�@              �?      *@              (@      �?      �?      �?                      �?     0r@      <@               @     0r@      :@     �p@      :@     �p@                      :@      8@             @T@            ���@    ���@    �z�@     ̔@     _�@     ȉ@     J�@     `�@     G�@      �@     �]@      �@              �@     �]@             Ѹ@              @      Z@              Z@      @             �@     �F@     ��@      C@     ��@               @      C@      �?      C@              C@      �?              �?             @c@      @      @      @      @                      @     `b@       @     �`@      �?     �`@                      �?      ,@      �?      (@      �?      (@                      �?       @             �K@     �@     �G@     �@      @      @               @      @      �?              �?      @             �E@     `@      5@     �d@             �d@      5@              6@     �t@             �t@      6@               @      �?              �?       @             p�@    �7�@     Pp@     �@      @      �?      @                      �?     p@      �@             ��@     p@       @      2@      �?      @              (@      �?      (@                      �?     �m@      �?     @\@      �?      S@      �?      S@                      �?     �B@             �_@             ̜@    ���@     @�@     ��@             ��@     @�@      ,@     �@              *@      ,@              ,@      *@             �A@     (�@             �@     �A@     @Q@               @     �A@     �N@             �L@     �A@      @      9@              $@      @      @      @      @                      @      @        �t�bubhhubehhub.