���'      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�K*�min_impurity_decrease�G        �min_impurity_split�N�class_weight�N�	ccp_alpha�G        �n_features_in_�K�n_features_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�h�scalar���h'C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h'�C       �t�bK��R�}�(h	K�
node_count�K�nodes�hhK ��h��R�(KK��h$�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hJh'K ��hKh'K��hLh'K��hMh$�f8�����R�(Kh(NNNJ����J����K t�bK��hNhXK ��hOh'K(��hPhXK0��uK8KKt�b�B�         H                  �th�?y�Q��?l�         ��A       5                 ����?�WS��?��         $"A                         �'��?��i��?�W         �_A                        ��� @b�)�7��?p4         ��A                        �?Z�?���BM��?�*         ��A       	                 0(*�?���_��?I          $�A                        ���?h~IZ���?�         �A������������������������       ���{��?�         �A������������������������       �D�1�J��?             7@
                        ��,�?��s���?K            �R@������������������������       �                     @������������������������       ��t�h���?E            @Q@                         n��?iG�����?�
           l�@                        �)d�?(�����?�
           b�@������������������������       �                     (@������������������������       ��%�t7��?�
           J�@������������������������       �                     @                        @��?H���j�?q	           �@                        ��?�@?��?R           H�@                        p�� @�>�<^ȷ?K           X�@������������������������       �|%��b�?             .@������������������������       �        <           ��@                         }ٚ����]���?           pp@������������������������       ����P#��?�            `j@������������������������       �vUb̙�?4             J@                        pEؿs��>I�?           |�@                        ��?�^��h�?P             T@������������������������       ���hX���?=            �N@������������������������       ��f1�a�?             3@                        PE� @�F�ոm�?�           <�@������������������������       ��Z���?
             $@������������������������       �X:dN�?�           �@!       ,                 @��?�.y;]��?u#          ���@"       '                 ��?��qa��?u           �@#       &                 `z��?�š?�           ��@$       %                 ���̿���s�?             :@������������������������       �                      @������������������������       �V�-���?             8@������������������������       �        �           l�@(       )                 ����?/['��U�?�           (�@������������������������       �                     @*       +                 `���?s��fl6�?�           ��@������������������������       ����Hi�?�            �a@������������������������       �f�(����?           ��@-       .                 `�y�x?����?             �@������������������������       �                      @/       2                 ��*Ϳ&.l«�?�           ��@0       1                 P&/Ϳ�X��P�?�            �j@������������������������       �̀M���?�             i@������������������������       ��n$����?             .@3       4                 zͿuS�U��?!           !�@������������������������       �T$?���?�             a@������������������������       �z	�[��?�           ��@6       7                 ��?x�����?�0           R�@������������������������       �        l#           ��@8       A                 0&a�?�.���?8           p�@9       :                 ` 3�?Ea�V�?�           ��@������������������������       �                     2@;       >                 ���%@p_Ǧc�?�           ��@<       =                 0u�@�
r�;o�?�           X�@������������������������       �U�u�e�?�           <�@������������������������       �������?             ,@?       @                  b&տ��S=�]�?             ;@������������������������       �                     (@������������������������       ��n$����?             .@B       C                 @��?$�A>���?_            �W@������������������������       �        '            �C@D       E                 �{�?̰����?8             L@������������������������       �                     @F       G                 `���?&[Z7��?4             J@������������������������       �                     @������������������������       �bD����?1            �H@I       d                 wؿ��ϧ��?�n          ���@J       [                 @��?�rg��?(           P�@K       L                 @��? ΢J�w�?�	           >�@������������������������       �        �            �l@M       T                 2��?ؓ���?�           p�@N       Q                 �vBɿ��`���?6           l�@O       P                 @�ٿ|��"��?�           H�@������������������������       ���Aޤ�?T           @u@������������������������       �l(�<��?u           ��@R       S                 ��	ؿ"���(e�?m           ��@������������������������       �w��6S�?h           ��@������������������������       �                     @U       X                 0��ٿ\�H�[�?�            @`@V       W                 Ш�ٿ������?             @������������������������       �|%��b�?             @������������������������       �                     @Y       Z                 �wJٿ�.� ���?{            �^@������������������������       �                     (@������������������������       ��t�W!�?o            �[@\       ]                 ��'@���3r�?�           H�@������������������������       �                   ��@^       _                 �L�?;�" E��?k            �Z@������������������������       �        Z            �V@`       c                 PrqؿB���-��?             1@a       b                 ���@JQe1���?             ,@������������������������       �.a�� �?             &@������������������������       �|%��b�?             @������������������������       �                     @e       n                 ���?ư�f���?�a          �n�@f       g                 ��� @6?UR��?yE          @^�@������������������������       �        �>          �s�@h       i                 `���?�����?�           H�@������������������������       �        &           ��@j       m                 ��?�,���?l           �v@k       l                 @_�@��nB���?\           �u@������������������������       �f�{4��?J           �t@������������������������       �|%��b�?             2@������������������������       �                     0@o       x                 @���?]&7uqo�?B           B�@p       q                 ��� @����e�?U           U�@������������������������       �        �           ��@r       u                 ��@�u׏\��?�            �f@s       t                 ��@���Z���?
             $@������������������������       �M�)9��?	             "@������������������������       �                     �?v       w                 �@_p�����?�            �e@������������������������       ��9>����?             <@������������������������       ��Y�Y��?�             b@y       ~                 ��?�<vmzd�?�           ��@z       }                 0'U-@�EzJ��?�           ��@{       |                 p+�%@#�Z����?�           ��@������������������������       �@��~X��?�           4�@������������������������       �� �2���?             9@������������������������       �                     @������������������������       �        C            �P@�t�b�values�hhK ��h��R�(KKKK��hX�B�      `��@    ��	A    T�@    @�A    P��@     XA    0��@    ��A    �7�@     �A    � �@    �A     ��@    ��A    ���@    @�A      @      4@      E@     �@@      @              B@     �@@     x�@     �@     P�@     �@              (@     P�@     �@      @             ��@     ȏ@     Ќ@      g@     �@      $@      @      $@     ��@             @V@     �e@     �S@     �`@      $@      E@     �}@     �@     �P@      ,@     �M@       @      @      (@     �y@     ��@       @       @     @y@     ��@     �@     �@     6�@     Ђ@     ��@      &@      .@      &@               @      .@      "@     l�@             `u@     x�@      @             �t@     x�@      A@      [@     �r@     0~@     \�@     R�@               @     \�@     B�@     @V@     �_@     �S@     �^@      &@      @     ��@     F�@      =@     �Z@     ��@     p�@     .�@     ��@     ��@             ��@     ��@     ؒ@     F�@              2@     ؒ@     "�@     Ȓ@     �@     ��@     ؟@      $@      @      @      7@              (@      @      &@      M@     �B@     �C@              3@     �B@      @              .@     �B@      @              (@     �B@     Ԗ@    �K�@     Ї@     \�@     ��@     ��@             �l@     ��@     �@     ��@     ��@     0s@     ��@      `@     `j@     @f@     0|@      z@     X�@     �y@     X�@      @              ?@     �X@      @       @      �?       @      @              :@     @X@              (@      :@     @U@      @     �@             ��@      @     @Y@             �V@      @      &@      @      &@      �?      $@       @      �?      @             ؅@     ��@     @`@    �=�@            �s�@     @`@     @�@             ��@     @`@     @m@     @`@     @k@     �]@     �j@      (@      @              0@     ȁ@     	�@     �O@     �@             ��@     �O@     �]@       @       @       @      �?              �?     �K@     @]@      @      8@     �I@     @W@     �@     ��@     �@     ��@     `@     ��@     0@     Ќ@      @      6@      @                     �P@�t�bub�_sklearn_version��0.24.2�ub.