���      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �min_impurity_split�N�class_weight�N�	ccp_alpha�G        �n_features_in_�K�n_features_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�h�scalar���h'C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h'�C       �t�bK��R�}�(h	K�
node_count�KC�nodes�hhK ��h��R�(KKC��h$�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hJh'K ��hKh'K��hLh'K��hMh$�f8�����R�(Kh(NNNJ����J����K t�bK��hNhXK ��hOh'K(��hPhXK0��uK8KKt�b�B�         "                  BHAhSVo�?l�         ��A                          �A��ǻv�?�t         P�A                         xA���?���?�:         ��A                         �wA  ����>�*         h�A������������������������       �        �*         L�A                         xA؇���X�?             @������������������������       �                     �?������������������������       �                     @	       
                    �?������?�           ¯@������������������������       �        ^           x�@                           �?
w����?�
           �@                           �?�g`�S��?�           x�@������������������������       �        (           ��@������������������������       �        �            �f@                          P��@0���[�?�           (�@                           �?��(�?q            @\@������������������������       �        d             Y@������������������������       �                     *@������������������������       �        4           ��@                           �?(M���r�?�9          ���@                           �?��ۖ��?�%          ���@                         �xA@�-	�?8           p�@������������������������       �                   �@                           �?r�q��?0             H@������������������������       �        (             D@������������������������       �                      @                           �?�}"�F�?�           ��@������������������������       �        %           %�@������������������������       �        \           ��@                         �xA�E�n4��?             �@������������������������       �        �           ٳ@        !                    �?@�j;��?G            �Q@������������������������       �        A            @P@������������������������       �                     @#       4                    �?�b�S���?؂           [�@$       1                   n�A����# �?�-          ���@%       ,                   �x�@|q
����?�+           ��@&       )                    �?d���r�?<           �@'       (                    �?���tT��?\           ��@������������������������       �        �           p�@������������������������       �        n            �[@*       +                  �hA �.�?Ƞ?�            ~@������������������������       �        �           �}@������������������������       �                      @-       .                  BxA@�X�
B�?�&           A�@������������������������       �        �%           ��@/       0                    �?���.�d�?�            �a@������������������������       �        �            �`@������������������������       �        	             "@2       3                    �?�c�Չ��?A           �@������������������������       �                   @�@������������������������       �        9            �L@5       6                    �?��&�=v�?�T          @6�@������������������������       �        CL          ��@7       >                   z�AP<B�v�?�           ,�@8       9                  :yA@��!�Q�?4           h�@������������������������       �                   ,�@:       ;                    �?�q�q�?             >@������������������������       �                     3@<       =                    �?�C��2(�?             &@������������������������       �                     �?������������������������       �        
             $@?       @                    �?j�Je���?b            �X@������������������������       �        A            @P@A       B                  �gA�FVQ&�?!            �@@������������������������       �                     ?@������������������������       �                      @�t�b�values�hhK ��h��R�(KKCKK��hX�B0      � A     ��@    �]A     �@    ��A     4�@    d�A      �?    L�A              @      �?              �?      @             ��@     0�@     x�@             ��@     0�@     �f@     ��@             ��@     �f@             �@      Y@      *@      Y@              Y@      *@             ��@            ���@     ��@     خ@     M�@      �@      D@     �@               @      D@              D@       @             ��@     %�@             %�@     ��@             ߳@     @P@     ٳ@              @     @P@             @P@      @            �]�@    @��@     >�@     �@    �!�@     ؋@     0�@     ��@     �[@     p�@             p�@     �[@             �}@       @     �}@                       @    ���@     �`@     ��@              "@     �`@             �`@      "@             �L@     @�@             @�@     �L@             ~�@    �&�@            ��@     ~�@     �U@     @�@      4@     ,�@              $@      4@              3@      $@      �?              �?      $@              ?@     �P@             @P@      ?@       @      ?@                       @�t�bub�_sklearn_version��0.24.2�ub.