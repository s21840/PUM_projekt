��      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�K*�min_impurity_decrease�G        �min_impurity_split�N�class_weight�N�	ccp_alpha�G        �n_features_in_�K�n_features_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�h�scalar���h'C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h'�C       �t�bK��R�}�(h	K�
node_count�K5�nodes�hhK ��h��R�(KK5��h$�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hJh'K ��hKh'K��hLh'K��hMh$�f8�����R�(Kh(NNNJ����J����K t�bK��hNhXK ��hOh'K(��hPhXK0��uK8KKt�b�B�                          ��¯?      �?��          ���@                         @���?�������?'�          ���@                        �p�?���e��?@m           P�@������������������������       �        �e          �r�@                        �@5�v��� ��?v           ؝@������������������������       �        �            @b@       
                 ���?n�b�Ef�?�           ��@       	                 
�_�?}S����?1           Ę@������������������������       �                    ��@������������������������       �                     1@                        <j<�^� ��?�            `f@������������������������       �        ^            �W@������������������������       �        U            @U@                        ���?��t�;�?�           �@                        �@5�@J9���?�           ��@                        ���?���N�\�?Y           �u@������������������������       �        .           �r@������������������������       �        +            �E@                        
�_�?�iR�ܹ?G           G�@������������������������       �        �           ��@������������������������       �        K            �R@                        �/��?I�9����?G           8�@������������������������       �                   �@������������������������       �        D             Q@       (                 �@5�7b��#,�?�V          ���@       !                  0��ۿ��{F�?C	           ��@                        ���?�*DQ���?           ��@                        
�_�?���8��?�           ��@������������������������       �        �           �@������������������������       �                     ,@                         ����?��%!��?/            �G@������������������������       �        '            �C@������������������������       �                      @"       %                  б��?�wMl�K�?$           ��@#       $                 ��?��6�?           d�@������������������������       �        �           ��@������������������������       �        �             `@&       '                 
�_�?��㛙�?           X�@������������������������       �                   @�@������������������������       �                     @)       *                 
�_�?ܪ����?DM           Q�@������������������������       �        'L          �	�@+       0                  �Ci�?�5@k��?           �q@,       -                 ���?�I>X���?�             j@������������������������       �        �             h@.       /                 �(u@�X)��?             0@������������������������       �                     .@������������������������       �                     �?1       2                 ���?���E�a�?L             S@������������������������       �        D             Q@3       4                 l}��?c�YB�d�?              @������������������������       �                     @������������������������       �                     �?�t�b�values�hhK ��h��R�(KK5KK��hX�BP      ���@    ���@    ���@     �@    ���@     ��@    �r�@              o@     ��@     @b@             �Y@     ��@      1@     ��@             ��@      1@             @U@     �W@             �W@     @U@             ��@     k�@     �w@     '�@     �r@     �E@     �r@                     �E@     �R@     ��@             ��@     �R@             �@      Q@     �@                      Q@     d�@    �{�@     ��@     ̕@     �J@     P�@      ,@     �@             �@      ,@             �C@       @     �C@                       @     ،@     H�@     ��@      `@     ��@                      `@      @     @�@             @�@      @              i@    ��@            �	�@      i@      U@     @h@      .@      h@              �?      .@              .@      �?              @     @Q@              Q@      @      �?      @                      �?�t�bub�_sklearn_version��0.24.2�ub.