���      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �min_impurity_split�N�class_weight�N�	ccp_alpha�G        �n_features_in_�K�n_features_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�h�scalar���h'C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h'�C       �t�bK��R�}�(h	K�
node_count�K-�nodes�hhK ��h��R�(KK-��h$�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hJh'K ��hKh'K��hLh'K��hMh$�f8�����R�(Kh(NNNJ����J����K t�bK��hNhXK ��hOh'K(��hPhXK0��uK8KKt�b�B�	                          �\�?      �?��          ���@       	                  �@��?�l���?)�           ��@                        �h��?	��|��?gm          �Y�@������������������������       �        �e          �{�@                        @��&���a��?x           ��@������������������������       �        �            �`@                        �W��?'�*�(<�?�           Л@������������������������       ��q�Q��?E           �@������������������������       �]EZ�%��?�            �e@
                        �W��?���m�#�?�           ¹@                        @����@p��?�           ��@                        �#��?*�s��t�?f           `v@������������������������       �        9           �s@������������������������       �        -            �F@                        ٍ�?!2���?,           ,�@������������������������       �        �           �@������������������������       �        A            @P@                        p�>�?X R&ڻ�?0           ��@������������������������       �        �           `@������������������������       �        :             M@       $                 @��$�3�) �?�V          @��@                         `�	ٿ��n�z;�?c	           Ƣ@                        �W��?RX�-��?"           �@                        ٍ�?dV
�?�           ��@������������������������       �        �           P�@������������������������       �                     (@                        @Ti�?�v*gjc�?,             F@������������������������       �        &             C@������������������������       �                     @       !                  ���?��1�Z]�?A           �@                         ���?(�Y$��?           d�@������������������������       �        �           �@������������������������       �        |             _@"       #                 ٍ�?�~t
&��?(           @�@������������������������       �                     �@������������������������       �                      @%       &                 ٍ�?bY�
�?"M          �H�@������������������������       �        L           �@'       *                  � ��?�Q�?           �p@(       )                 �k��?��~���?�            �h@������������������������       �        �            �f@������������������������       ��X)��?             0@+       ,                 �W��?��W�I��?G            �Q@������������������������       �        A            @P@������������������������       �                     @�t�b�values�hhK ��h��R�(KK-KK��hX�B�      ���@    ���@    ���@     �@    ���@     T�@    �{�@             `l@     T�@     �`@             �W@     T�@      0@     Ԙ@     �S@      X@     ��@     R�@     �w@     �@     �s@     �F@     �s@                     �F@     @P@     �@             �@     @P@             `@      M@     `@                      M@     T�@     |�@     ��@     0�@      I@     ��@      (@     P�@             P�@      (@              C@      @      C@                      @     (�@     ��@     �@      _@     �@                      _@       @      �@              �@       @             �g@     �@             �@     �g@      T@      g@      .@     �f@              �?      .@      @     @P@             @P@      @        �t�bub�_sklearn_version��0.24.2�ub.