��     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �min_impurity_split�N�class_weight�N�	ccp_alpha�G        �_sklearn_version��0.24.2�ub�n_estimators�K�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK�verbose�K �
warm_start��hN�max_samples�NhhhKhKhKhG        h�auto�hNhG        hNhG        �n_features_in_�K�n_features_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h-�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhKhKhKhG        hh%hNhJc��8hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��h6�f8�����R�(Kh:NNNJ����J����K t�b�C              �?�t�bh>h*�scalar���h9C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hK�
node_count�K��nodes�h,h/K ��h1��R�(KK���h6�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hkh9K ��hlh9K��hmh9K��hnhJK��hohJK ��hph9K(��hqhJK0��uK8KKt�b�BX)         @                 ����bˢ��?�           ��@       7                  �;0�?�Ϝ�K-�?i           ��@       $                 @���?p?t�P�?<           ��@       #                  ��?�d��D��?�           �@                        0���?���-��?a           �@������������������������       �        &           0}@       "                 @��?���;+"�?;            �S@                         � �?��(@��?4            �Q@	                        �T�?Fx$(�?"             I@
                          g�ٿ�n_Y�K�?             *@������������������������       �                     @������������������������       �                      @                        `@��?V������?            �B@������������������������       �        
             *@                        �[X�?r�q��?             8@                          q�ڿ      �?              @������������������������       �                      @������������������������       �                     @                        ���?     ��?             0@������������������������       �                     @                        ps�?�q�q�?             (@������������������������       �z�G�z�?             @������������������������       �؇���X�?             @                        �=�?�z�G��?             4@������������������������       �                     @                         �X�?���Q��?             .@������������������������       �                     �?                        �2��?X�Cc�?             ,@������������������������       �                      @                        p�@�?�q�q�?             (@������������������������       �                      @        !                 ����?�z�G��?
             $@������������������������       �                     @������������������������       �և���X�?             @������������������������       �                     "@������������������������       �        (            �O@%       &                  ��?�=ѱ?�            Pq@������������������������       �        �             m@'       6                  �KM˿�<ݚ�?            �F@(       5                  ��/Կ��}*_��?             ;@)       *                 `�7�?�q�q�?             8@������������������������       �                      @+       4                 ����?�GN�z�?             6@,       3                 ���?     ��?             0@-       2                  @!ڿd}h���?             ,@.       /                 �
�?      �?              @������������������������       �                      @0       1                  � vڿ      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �        
             2@8       ?                 �l2��B� ��?-            �Q@9       :                 �̀�@4և���?             E@������������������������       �                     <@;       <                  ��W�?d}h���?
             ,@������������������������       �                     $@=       >                 @���?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     <@A       �                 ��;�?B�h&��?N	           �@B       �                  ��?�P.^��?R           0�@C       �                  �0��?�k�Z��?�           �@D       c                 07�dIx���?�           l�@E       b                 ���l�G��=�?C            �^@F       K                 p1�迺�A���?B             ^@G       J                 �鿀��7�?             6@H       I                 ����q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     3@L       M                  �y�ۿJm_!'1�?3            �X@������������������������       �                      @N       W                  p��ٿr�q��?2             X@O       T                 @ט� �o_��?             9@P       Q                  Х�ڿ����X�?             @������������������������       �                     @R       S                  �3ڿ      �?             @������������������������       �                      @������������������������       �                      @U       V                 �d������H�?	             2@������������������������       �                     0@������������������������       �                      @X       ]                  @Iտ��UV�?&            �Q@Y       \                 `3p�h�����?             <@Z       [                  �=�ؿ      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     4@^       _                 �к�&^�)b�?            �E@������������������������       �                      @`       a                   �ѿ�p ��?            �D@������������������������       ��	j*D�?             *@������������������������       �@4և���?             <@������������������������       �                      @d       �                  p�bڿ wVX(6�?d           ��@e       �                  ��mڿ�p ��?|            �i@f       w                 Ўhۿ������?u            @h@g       t                 ��
ݿ�� =[�?S             a@h       m                  �0YۿX�GP>��?O            �_@i       j                 ���߿�&=�w��?            �J@������������������������       �                     G@k       l                  ��ۿ����X�?             @������������������������       �                      @������������������������       �                     @n       q                 @���?��A��?4            �R@o       p                  �S=ۿ4��?�?$             J@������������������������       �                     �?������������������������       ��:�]��?#            �I@r       s                   d�ڿ���|���?             6@������������������������       �      �?             0@������������������������       �                     @u       v                  ���ڿ�<ݚ�?             "@������������������������       �                     @������������������������       �                      @x       {                  ��xۿXB���?"             M@y       z                  �ӑۿ      �?             @������������������������       �                     @������������������������       �                     �?|                         `n�ڿ@3����?              K@}       ~                  ��ڿ�nkK�?             7@������������������������       �                     6@������������������������       �                     �?������������������������       �                     ?@�       �                  �,kڿ�eP*L��?             &@������������������������       �                     @�       �                 h6Vٿ      �?              @�       �                  иeڿr�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                 0@����q"���?�           P�@�       �                  PɁտ�S�L��?�           ��@�       �                 @���?4��?�?O           @�@�       �                 �I�俄YM_b�?�            �w@�       �                   /�ٿ@���|N�?L             `@�       �                 p��R���Q�?             4@������������������������       �                     "@������������������������       ����!pc�?             &@�       �                 Jk�HQ˄�ľ?@            @[@������������������������       �                     ;@������������������������       �ĴF���?0            �T@�       �                 ���T���RB�?�             o@������������������������       �                     @�       �                  @T�տ 4�"=[�?�            �n@������������������������       ���2(&�?�            @n@������������������������       �                     @������������������������       �        b            �a@�       �                 ��b��=QcG��?�           �@�       �                 @��p�
��ѻ?�           ��@�       �                  @@��?xP�Fֺ�?5            @V@�       �                 @���?�Ra����?4             V@������������������������       �д>��C�?!             M@������������������������       �                     >@������������������������       �                     �?�       �                 @���?�-@�w��?K           0�@�       �                  0<$�?��r��?�            pv@������������������������       �؇D^��?�            �t@������������������������       ��חF�P�?             ?@������������������������       �        a            �c@������������������������       �                     @������������������������       �                    �D@�       �                 �^t��.��?Q           H�@�       �                  |��j��b�?'            �M@�       �                 @���?�h����?&             L@������������������������       �        $            �J@������������������������       �                     @������������������������       �                     @�       �                 @���? ��WV�?*           �~@������������������������       �                   �}@������������������������       �                     3@������������������������       �        Z            �b@�       �                 P@�*@@��� ��?�           ��@�       �                  ��? C��»�?�           ��@������������������������       �        �           h�@�       �                 @���?z�G�z�?             .@�       �                  �g�ڿ�θ�?	             *@������������������������       �                     �?�       �                  ���?r�q��?             (@�       �                 P�'�?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�t�b�values�h,h/K ��h1��R�(KK�KK��hJ�B�       �@     ��@     (�@     �U@     ��@      L@     ��@      G@     @@      G@     0}@             �@@      G@     �@@     �B@      3@      ?@       @      @              @       @              &@      :@              *@      &@      *@      @       @               @      @              @      &@              @      @      @      @      �?      �?      @      ,@      @      @              "@      @              �?      "@      @       @              @      @               @      @      @      @              @      @              "@     �O@             �p@      $@      m@             �A@      $@      1@      $@      1@      @               @      1@      @      &@      @      &@      @      @      @       @              @      @      @                      @      @                       @      @                      @      2@             �C@      ?@     �C@      @      <@              &@      @      $@              �?      @              @      �?                      <@     ,�@     �@     �@     ��@     ��@     ��@     <�@     �a@     @Y@      5@     @Y@      3@      5@      �?       @      �?       @                      �?      3@              T@      2@               @      T@      0@      2@      @       @      @              @       @       @       @                       @      0@       @      0@                       @      O@      "@      ;@      �?      @      �?              �?      @              4@             �A@       @               @     �A@      @      "@      @      :@       @               @     ��@     �]@     �e@      >@     @e@      8@     �\@      6@      \@      .@     �I@       @      G@              @       @               @      @             �N@      *@     �G@      @              �?     �G@      @      ,@       @       @       @      @               @      @              @       @              L@       @      @      �?      @                      �?     �J@      �?      6@      �?      6@                      �?      ?@              @      @              @      @      @      @      �?      @                      �?               @     �@     @V@     H�@     @V@     `}@      I@     �t@      I@     �]@      $@      1@      @      "@               @      @     �Y@      @      ;@             �R@      @      j@      D@              @      j@     �B@      j@     �@@              @     �a@             ��@     �C@     ��@     �A@     �S@      &@     �S@      $@      H@      $@      >@                      �?     �~@      8@     �t@      8@     Ps@      3@      :@      @     �c@                      @     �D@              9@     ��@      @     �J@      @     �J@             �J@      @              @              3@     �}@             �}@      3@             �b@              .@     t�@      (@     t�@             h�@      (@      @      $@      @              �?      $@       @      $@      �?      $@                      �?              �?       @              @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh%hNhJ�H hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK˅�hi�Bh,         �                 ���?      �?           ��@                        ����joq�M�?n           J�@                        @���? o6��%?           ��@                        p�h��O"9��?a           ��@������������������������       �        �            Ps@                         `�~	@`׀�:M�?�            �k@                         ��W�?�������?�            �k@������������������������       �        �             k@	       
                  �Wa@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        �            �o@                         �0��?l�D���?l           &�@       :                   bֿ��.A��?           ę@                        б����&�?�           ��@                        ���      �?             @������������������������       �                     �?������������������������       �                     @       +                 @���? ��#��?�           p�@       *                  N�@�"�t�(�?e           p�@       )                  �ycֿ��̃��?]           ��@                          `�uڿ�m�F�?[           �@                        P������a�n`�?c            `c@                        `@�㿈˹�m��?b             c@                        ��~�0�,���?,            �P@������������������������       �      �?             0@������������������������       ����J��?!            �I@                         ��?�t����?6            @U@������������������������       �d1<+�C�?-            @R@������������������������       �        	             (@������������������������       �                     @!       "                  �,kڿ8�v�l�?�             x@������������������������       �                     @#       &                  pL�ٿ��	W��?�            �w@$       %                  �,.ڿ�q��/��?6             W@������������������������       ��㙢�c�?             G@������������������������       ��nkK�?             G@'       (                  0h�ٿ�:7]4D�?�            r@������������������������       �                     @������������������������       �L���˚�?�            �q@������������������������       �                      @������������������������       �                     .@,       3                 P���Cc}�?�             l@-       0                 �����q�q�?             8@.       /                  �EUۿ@�0�!��?	             1@������������������������       �                     @������������������������       �                     ,@1       2                  �G�ڿ����X�?             @������������������������       �                     @������������������������       �                      @4       9                  ��?�c�ZB�?�             i@5       8                  �ܩڿ�b��fl�?z             g@6       7                  �6�ڿ�#-���?            �A@������������������������       �                     @@������������������������       �                     @������������������������       �        ^            �b@������������������������       �                     0@;       ~                 @���?hx�,���?           ��@<       K                 �}&�f�\�~�?]           ��@=       F                 @Z6迊c�Α�?             =@>       E                  ��?�LQ�1	�?             7@?       @                  ��Hѿ��2(&�?             6@������������������������       �                      @A       D                 @R��P���Q�?             4@B       C                 �=��z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             .@������������������������       �                     �?G       H                  �Ͽr�q��?             @������������������������       �                     @I       J                  �,��q�q�?             @������������������������       �                      @������������������������       �                     �?L       g                  �3׿�s#}c�?K           ��@M       X                 �Z��=QcG��?           pz@N       W                 ���濸��H��?3             U@O       R                  ���տ��Lɿ��?2            �T@P       Q                  ��/ֿ�q�q�?             @������������������������       �                     �?������������������������       �                      @S       V                  ��?p=
ףp�?0             T@T       U                 ���pH����?)            �P@������������������������       �85�}C�?$            �N@������������������������       ��q�q�?             @������������������������       �                     *@������������������������       �                     �?Y       f                  ��?@��Pc�?�            0u@Z       a                  �RԿ�&����?�            `s@[       ^                  p�)Կ�:pΈ��?"             I@\       ]                 @	�ῴC��2(�?             F@������������������������       �Pa�	�?            �@@������������������������       ����!pc�?             &@_       `                 p��      �?             @������������������������       �      �?             @������������������������       �                      @b       c                 ��T� ��WV�?�            @p@������������������������       �        >            �W@d       e                  ����� ,U,?��?h            �d@������������������������       ��v�ɱ?B            �[@������������������������       �lGts��?&            �K@������������������������       �                     =@h       o                  �<sͿ��#:���?=            �[@i       j                 `��ֿ@4և���?             E@������������������������       �                      @k       n                  PɁտ�(\����?             D@l       m                  pg�տr�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     A@p       w                 y�ӿH�V�e��?"             Q@q       r                 ���Կ��S���?             .@������������������������       �                     @s       t                   c/ƿz�G�z�?             $@������������������������       �                     @u       v                  x�`���q�q�?             @������������������������       �                      @������������������������       �                     @x       y                 �Brɿ���C��?            �J@������������������������       �                     :@z       {                 0��ȿ�<ݚ�?             ;@������������������������       �                     �?|       }                 p�ѭ����B���?             :@������������������������       ������H�?             2@������������������������       �      �?              @������������������������       �        �            �r@�       �                  ��?y����?e           �@�       �                 �؍?�f�����?^           Ȁ@�       �                 ��㿸w�>τ�?X           p�@�       �                 @���?0�K炇�?�            pp@������������������������       �        �             p@������������������������       �                     @�       �                 �x}��Qɕ9��?�            pp@������������������������       �                      @�       �                 @���?�D�
Q;�?�            Pp@������������������������       �        �             o@������������������������       �        	             *@�       �                 ����?���!pc�?             &@������������������������       �                     @������������������������       �                      @������������������������       �                     "@�       �                 ���濘�{Oӷ?�           l�@�       �                  �ڿ"�����?~            �i@�       �                  ��?�}�+r��?0             S@�       �                 @���?`2U0*��?/            �R@������������������������       �        ,            �Q@�       �                  `:Tۿ���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                  ��?-"� ��?N            ``@�       �                 ����?v�\!L^�?I            @^@�       �                 @���?���y4F�?             3@�       �                 @�=�?      �?             (@�       �                 ��_�?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                  ���ؿ؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                 p�P�?��.k���?=            �Y@�       �                 `���?�lg����?            �E@������������������������       �                     @�       �                  ���?D�n�3�?             C@�       �                  0ġٿ���!pc�?             6@�       �                 0| �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                 �I��?r�q��?
             2@�       �                 @���?�z�G��?             $@�       �                  ^zͿ      �?              @������������������������       �                     @������������������������       �      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     0@�       �                   f��?:���W�?%            �M@�       �                 @���?�����?             E@�       �                 0f<�?H%u��?             9@������������������������       �                     5@�       �                  ��)׿      �?             @������������������������       �                     �?������������������������       �                     @�       �                  (�ѿ�IєX�?             1@������������������������       �                     (@�       �                  �KM˿z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     1@������������������������       �                     $@�       �                 ��'@ 4��`~?           0�@�       �                 �ҳ�?�>y~�Xy?           ,�@�       �                  ��?@��� ��?e            �@������������������������       �        _           ��@�       �                 @�?r�q��?             @������������������������       �                     @�       �                 �W�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        �           ��@������������������������       �                     �?�t�bh~h,h/K ��h1��R�(KK�KK��hJ�B�       ��@     ��@     �@     ��@     x�@      @     ��@      @     Ps@             `k@      @     `k@      �?      k@               @      �?              �?       @                       @     �o@             ��@     ؄@     X�@     `c@     X�@     �Y@      �?      @      �?                      @     P�@      Y@     P}@     @V@     `|@     @V@     `|@     �U@     �a@      .@     �a@      (@     @P@       @      .@      �?      I@      �?     �R@      $@     �O@      $@      (@                      @     �s@      R@              @     �s@     �P@     �T@      $@      C@       @      F@       @      m@     �L@              @      m@      K@               @      .@             �j@      &@      0@       @      ,@      @              @      ,@               @      @              @       @             �h@      @     �f@      @      @@      @      @@                      @     �b@              0@             X�@      J@     �@      J@      5@       @      4@      @      3@      @               @      3@      �?      @      �?      @                      �?      .@              �?              �?      @              @      �?       @               @      �?             �~@      F@     �x@      ;@     �R@      $@     �R@      "@      �?       @      �?                       @     @R@      @      N@      @      L@      @      @       @      *@                      �?      t@      1@     Pr@      1@     �E@      @      D@      @      @@      �?       @      @      @      @      @      �?               @     @o@      $@     �W@             �c@      $@     �Z@      @     �H@      @      =@             @W@      1@     �C@      @               @     �C@      �?      @      �?      @                      �?      A@              K@      ,@      @       @      @               @       @              @       @      @       @                      @     �G@      @      :@              5@      @              �?      5@      @      0@       @      @      @     �r@              A@      �@      9@      �@      6@     �@      @      p@              p@      @              .@      o@       @              *@      o@              o@      *@              @       @      @                       @      "@             @V@     �@     �T@      _@      @      R@      @      R@             �Q@      @       @               @      @              �?             �S@      J@     @Q@      J@      .@      @      "@      @      @      @      @                      @      @              @      �?              �?      @              K@      H@      0@      ;@              @      0@      6@      0@      @      �?      @              @      �?              .@      @      @      @      @      @      @              �?      @       @               @                      0@      C@      5@      C@      @      6@      @      5@              �?      @      �?                      @      0@      �?      (@              @      �?              �?      @                      1@      $@              @     �@      @     �@      @     ��@             ��@      @      �?      @               @      �?              �?       @                     ��@      �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh%hNhJ�O�^hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK�hi�B(5         R                 ����r�q��?�           ��@       7                 @���?x�ۈp�?�           �@       "                  �.�ڿ؇���X�?�           P�@       	                  0Áۿ�U���?K             _@                          ��ۿ8�Z$���?
             *@                        pw��?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     "@
       !                  ��?^H���+�?A            �[@                         Ћۿy�w[��?@            @[@                        ��E��.��<�?%            �P@������������������������       �                     1@������������������������       �                     I@                         �M�ڿ�G��l��?             E@                        `󁱿@�0�!��?             1@������������������������       �                     ,@������������������������       �                     @                         ���ڿ�+e�X�?             9@                         �H�ڿףp=
�?             $@                         ���ڿz�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                         ���ڿ�q�q�?	             .@                         �z�ڿ�q�q�?             @                         ���?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                          �i�������H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                      @#       6                  ��?���)%�?o           p�@$       +                 0���?@?i����?G           P�@%       *                  0mp@ UGH�?!           `}@&       '                  ���?�&���q?           0}@������������������������       �                   �|@(       )                  @���?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @,       5                   f��?��
ц��?&             J@-       .                  �0�˿��S�ۿ?             >@������������������������       �                     3@/       4                  �Ɵ��"pc�
�?
             &@0       1                  `)�ſ�q�q�?             @������������������������       �                     �?2       3                 �I��?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     6@������������������������       �        (             Q@8       M                  P�N�?0G���ջ?�            �s@9       <                  p`�ۿ�Ń��̧?�            `r@:       ;                  `қۿ      �?             @������������������������       �                     @������������������������       �                     �?=       >                 `��?@��t��?�             r@������������������������       �        �            �n@?       L                  ��?�r����?!            �F@@       K                  �KM˿؇���X�?             E@A       J                  p1�ҿ�θ�?             :@B       C                 ����?r�q��?             8@������������������������       �                      @D       I                  @!ڿ�C��2(�?             6@E       H                 �v�?����X�?             @F       G                 �
�?      �?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                     .@������������������������       �                      @������������������������       �        
             0@������������������������       �                     @N       Q                  ��t@b�2�tk�?             2@O       P                 ���ÿ     ��?             0@������������������������       �                     @������������������������       �                     &@������������������������       �                      @S       �                  ��?d2ҟp��?@	           |�@T       �                  �!��?=� ��?�           �@U       �                 ����?���g��?b           z�@V       �                 @���?����Ԅ�?�           (�@W       z                  �2�տ�g�ځ��?�           $�@X       e                  `�uڿRe�*��?]           h�@Y       d                 P���������?W            �b@Z       c                  ���ڿ�1h�'��?V            `b@[       b                  �J�ڿ��|���?7             V@\       _                  �I�ۿ �Cc}�?5             U@]       ^                 pI�      �?              @������������������������       �                     �?������������������������       �                     �?`       a                 @���������?3            �T@������������������������       �                     ?@������������������������       �>a�����?            �I@������������������������       �                     @������������������������       �                    �M@������������������������       �                     �?f       y                 `tÿ�)�ӯ��?           �y@g       l                  �,kڿ��r��?�            �w@h       k                  ��mڿz�G�z�?             @i       j                 Pc�      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @m       t                 @�(˿F2�y��?�            `w@n       q                  �����wy���?�             w@o       p                 ���      �?              @������������������������       �                     @������������������������       �                     @r       s                 @��z�G�z�?�            �v@������������������������       �        
             .@������������������������       �6@��]#�?�            �u@u       x                  �Xſ�q�q�?             @v       w                  �7ٿ      �?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                      @������������������������       �                     >@{       �                  ��h�?POͳF��?3           �}@|       �                 ���~���?           �y@}       �                 �s�L<8)��?�            �o@~       �                  `Rѿ�J�4�?6            �R@       �                  ��	Կ��R[s�?            �A@�       �                  ��*տ�IєX�?	             1@������������������������       ��q�q�?             @������������������������       �                     ,@�       �                 �}&�X�<ݚ�?             2@������������������������       �                     @������������������������       �����X�?             ,@�       �                 �s2���(\���?"             D@�       �                  @�|��      �?             @@������������������������       �                     :@������������������������       �r�q��?             @�       �                 �I�      �?              @������������������������       �                     �?������������������������       �؇���X�?             @�       �                 P�O忐��!5��?n            `f@�       �                 �wc�0G���ջ?             J@�       �                  @N�Կp���?             I@������������������������       �                     �?������������������������       �                    �H@������������������������       �                      @�       �                 ���U���?Q            �_@�       �                 �����Μ�5�?E            �[@������������������������       �(;L]n�?%             N@������������������������       �                     �I@�       �                 0o��      �?             0@������������������������       �                     �?������������������������       �                     .@�       �                 `��࿘�q縬�?g            �c@�       �                  ��ӿX�<ݚ�?             2@�       �                 ��؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                  �\ſ"pc�
�?             &@�       �                  Аʿ����X�?             @������������������������       �r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                  ��ѿ�{"z;m�?\            �a@�       �                 ���׿@3����?$             K@������������������������       �                     =@�       �                  `[�ҿ`2U0*��?             9@������������������������       ��8��8��?	             (@������������������������       �                     *@�       �                 ��ڿ\-��p�?8            �U@������������������������       �                    �@@�       �                  �~Wп�<ݚ�?'             K@������������������������       �                     @������������������������       �@�0�!��?&            �I@�       �                  ����?d�;lr�?(            �O@������������������������       �                     @�       �                 '��ܷ��?��?&             M@�       �                  Ў��?     ��?
             0@�       �                  �K��?@4և���?	             ,@������������������������       �                     @�       �                  ��?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                  ����?@4և���?             E@�       �                  �9��?d}h���?             ,@������������������������       �                     $@�       �                 H�ѿ      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     <@�       �                 0�翐�4J;�?           |@�       �                  ��ۿPN��T'�?             ;@�       �                 ���z�G�z�?             @�       �                 �R4�      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     6@�       �                  �}�ڿ@�'�W��?
           `z@�       �                 �J��8��8���?$             H@�       �                  ��]ۿ     ��?             0@������������������������       �                     @�       �                 �F��      �?             $@�       �                 �>��r�q��?             @�       �                  �G�ڿ�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @@������������������������       �        �            `w@������������������������       �        �           ̗@�       �                 ��⿰�ܲe6�?p           h�@�       �                  p�@�i��Lg�?�            pr@�       �                 ���� E��ۛ?�             r@�       �                 @���?���N8�?8             U@������������������������       �        5             T@������������������������       �                     @������������������������       �        y            �i@�       �                 @���?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                 @���?`<���?�            `r@������������������������       �        �             p@�       �                 p~Ү?�s��:��?             C@������������������������       �                     1@������������������������       �                     5@�       �                 `mO�?��r�#�?n            �f@�       �                 @���?�������?g            �d@�       �                 �H��? ��+&ɐ?K            @^@������������������������       �        I            �]@�       �                 ���?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                    �F@�       �                 @���?և���X�?             ,@�       �                  �؍�?���Q��?             $@�       �                 P�'�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh~h,h/K ��h1��R�(KK�KK��hJ�B0       �@     ��@     P�@      ^@      �@     �Y@      I@     �R@      &@       @       @       @       @                       @      "@             �C@      R@     �B@      R@      1@      I@      1@                      I@      4@      6@      ,@      @      ,@                      @      @      3@      �?      "@      �?      @              @      �?                      @      @      $@      @       @      �?       @      �?                       @      @              �?       @      �?                       @       @             ��@      <@     �~@      <@      }@      @      }@      �?     �|@              @      �?              �?      @                      @      <@      8@      <@       @      3@              "@       @      �?       @              �?      �?      �?              �?      �?               @                      6@      Q@             `r@      2@     �q@      @      @      �?      @                      �?     �q@      @     �n@             �C@      @      B@      @      4@      @      4@      @               @      4@       @      @       @       @       @      �?              �?       @      @              .@                       @      0@              @              @      &@      @      &@      @                      &@       @             ��@     ��@     �@     ��@     ��@     H�@     ��@     �c@     ��@     �b@     �|@     �X@     �`@      ,@     �`@      *@     �R@      *@     �R@      "@      �?      �?      �?                      �?     �R@       @      ?@             �E@       @              @     �M@                      �?     Pt@      U@     pr@      U@      �?      @      �?      �?              �?      �?                      @     `r@      T@     @r@      S@      @      @      @                      @      r@      R@      .@             q@      R@       @      @       @       @              �?       @      �?               @      >@             �z@      J@     @w@     �D@     �m@      2@     �O@      (@      :@      "@      0@      �?       @      �?      ,@              $@       @              @      $@      @     �B@      @      ?@      �?      :@              @      �?      @       @              �?      @      �?     �e@      @     �H@      @     �H@      �?              �?     �H@                       @      _@      @     @[@       @      M@       @     �I@              .@      �?              �?      .@              a@      7@       @      $@      @      �?              �?      @               @      "@       @      @      �?      @      �?                      @      `@      *@     �J@      �?      =@              8@      �?      &@      �?      *@             �R@      (@     �@@              E@      (@              @      E@      "@      J@      &@              @      J@      @      *@      @      *@      �?      @              @      �?              �?      @                       @     �C@      @      &@      @      $@              �?      @              @      �?              <@             �{@      "@      7@      @      �?      @      �?      �?              �?      �?                      @      6@             z@      @     �E@      @      &@      @      @              @      @      @      �?       @      �?              �?       @              @                      @      @@             `w@                     ̗@      7@     ��@      @     r@      @     �q@      @      T@              T@      @                     �i@       @      @              @       @              1@     Pq@              p@      1@      5@      1@                      5@     �e@      @     �d@      �?      ^@      �?     �]@               @      �?              �?       @             �F@               @      @      @      @      @      �?      @                      �?              @      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh%hNhJ���ThG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B�!         6                 ����JY�8���?�           ��@                         @��ڿ�����o�?           �@       
                  ��?���ȫ�?e            �d@                        @���?�z�Ga�?b             d@                        �Ҳ?���N��?D             ]@������������������������       �                    �K@������������������������       �        %            �N@       	                 ����?`���i��?             F@������������������������       �                    �E@������������������������       �                     �?������������������������       �                     @       5                  ��?0�#�	)�?           �@       "                 @���?���Ժ?�           8�@                        @p��?p�eU}�?F           �@                         0mp@@���a��?#           �|@                         p���?��ꤘ�?"           �|@������������������������       �                   �{@                          ��?@�0�!��?             1@������������������������       �                     �?                         ���?      �?             0@������������������������       �                     @                         @���?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @������������������������       �                     �?       !                  �0�?\�����?#            �K@                          �Q�?<���D�?            �@@                         PU���`Jj��?             ?@������������������������       �                     5@                        ���?z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �        
             6@#       ,                  �;0�?P���Q�?�            @p@$       %                 (��? Df@��?�             o@������������������������       �        �            �k@&       '                  �q�?d}h���?             <@������������������������       �                     @(       +                 E��?�nkK�?             7@)       *                 ���?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     3@-       4                   ��@���|���?             &@.       /                  ��g�?�<ݚ�?             "@������������������������       �                     @0       3                  ���?�q�q�?             @1       2                 ���?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �        1            �V@7       �                 ���?h�Nɪ��?V	           t�@8       s                 @���?�X3`!�?V           �@9       f                 ��л��$NL_�?$           0�@:       a                  ��¿�ŇR���?�           ��@;       ^                  �RO�?MZqi�?�           T�@<       ]                  ��?(� �!��?�           ��@=       T                 �v�ʿ�	CO���?n           ��@>       G                  pq�ҿԀHM���?[           ȍ@?       F                  ���ҿ�اt?�?�           x�@@       C                 �g3ؿ& nF�?�           h�@A       B                 �T,ٿh�+���?d           X�@������������������������       ���?�?]           ��@������������������������       ���
ц��?             *@D       E                  а ؿ�FVQ&�?-            �P@������������������������       ��KM�]�?             C@������������������������       �                     <@������������������������       �                      @H       M                  �������S�ۿ?�            �t@I       L                 �Y+�0m��5!�?o            �f@J       K                  Pi̿������?2            �T@������������������������       ��>����?             K@������������������������       �                     <@������������������������       �        =            �X@N       Q                  �⳽�p�"�0�?Z            �b@O       P                 �#��q�q�?             "@������������������������       �                      @������������������������       �؇���X�?             @R       S                  @[ر��#-���?T            �a@������������������������       �@�0�!��?             1@������������������������       ���p\�?H            �^@U       V                 @�ʿX�Cc�?             <@������������������������       �                     @W       \                  ���¿"pc�
�?             6@X       [                  ��Ŀ      �?             0@Y       Z                 @�Sǿz�G�z�?             .@������������������������       ����Q��?             @������������������������       �ףp=
�?             $@������������������������       �                     �?������������������������       �                     @������������������������       �        8             V@_       `                  ��?&_���?7           �~@������������������������       �        2           �}@������������������������       �                     .@b       e                  ���?�LQ�1	�?             7@c       d                 �-���և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     0@g       r                  ��?      �?;             X@h       q                  ����?���!pc�?5             V@i       j                 P����Pa�	�?*            �P@������������������������       �                     <@k       l                 �Z(���}�+r��?             C@������������������������       �                     �?m       p                 P�-���?�|�?            �B@n       o                 P=����8��8��?
             (@������������������������       �        	             &@������������������������       �                     �?������������������������       �                     9@������������������������       �                     6@������������������������       �                      @t       �                 @��޿`�E���?2           P~@u       �                  ��?���j�?�            @s@v       �                 ��߿��K˱F�?�            �q@w       ~                 �/���/R���?�            �q@x       y                  �*�ڿ@4և���?             E@������������������������       �                      @z       }                  `��ڿ�(\����?             D@{       |                  P��ڿ      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     B@       �                 �%+� B&���?�             n@�       �                  �}�ڿ@|����?�             m@�       �                 �J��ܷ��?��?             =@�       �                 �u���θ�?             *@�       �                  ��]ۿ�C��2(�?             &@������������������������       �                     @������������������������       �      �?             @������������������������       �                      @������������������������       �                     0@������������������������       �        �            �i@�       �                 ���      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     6@������������������������       �        l             f@�       �                  ��?���R�?            $�@������������������������       �        �           ؘ@�       �                 @���?p�ݯ��?             3@�       �                  <��?�q�q�?	             (@�       �                 �G�?����X�?             @�       �                 �W�?r�q��?             @�       �                 �B=�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh~h,h/K ��h1��R�(KK�KK��hJ�B�	       �@     r�@     �@     @Z@     �Y@      O@     �X@      O@     �K@     �N@     �K@                     �N@     �E@      �?     �E@                      �?      @             ��@     �E@     ��@     �E@     P~@      >@     �|@      @     �|@      @     �{@              ,@      @              �?      ,@       @      @              @       @               @      @                      �?      =@      :@      =@      @      =@       @      5@               @       @               @       @                       @              6@     �n@      *@     `n@      @     �k@              6@      @              @      6@      �?      @      �?      @                      �?      3@              @      @       @      @              @       @      @       @      �?       @                      �?              @       @             �V@             ��@     ��@     x�@     ��@     �@     H�@     ؍@     ��@     ��@     �@     H�@     �`@     ��@     �`@     ��@     �^@     X�@      Y@     X�@     �X@     �|@     �W@     p|@     �U@      @      @      O@      @      A@      @      <@                       @     @s@      6@      f@      @     �S@      @      I@      @      <@             �X@             ``@      2@      @      @       @              �?      @      `@      (@      ,@      @     �\@      "@      2@      $@              @      2@      @      (@      @      (@      @      @       @      "@      �?              �?      @              V@              .@     �}@             �}@      .@              @      4@      @      @              @      @                      0@      R@      8@      P@      8@      P@       @      <@              B@       @              �?      B@      �?      &@      �?      &@                      �?      9@                      6@       @             �}@      $@     �r@      $@     @q@      $@     @q@      @     �C@      @               @     �C@      �?      @      �?      @                      �?      B@             �m@      @     �l@      @      :@      @      $@      @      $@      �?      @              @      �?               @      0@             �i@              @      �?              �?      @                      @      6@              f@              (@     ��@             ؘ@      (@      @      @      @      @       @      @      �?       @      �?       @                      �?      @                      �?              @      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh%hNhJ��4hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK�hbh,h/K ��h1��R�(KK���hi�B8#         L                 ����u�ҕ��?�           ��@       	                  ��ڿ0�� �?�            �@                        �0��?�ՙ/�?b            `b@������������������������       �        :            �U@                        @���?��S�ۿ?(             N@                         ��?0�)AU��?&            �L@������������������������       �        %             L@������������������������       �                     �?������������������������       �                     @
       5                 @���? ��26��?;           ��@       *                  pQ�?xt��ʻ?�           ��@                        ���?PaRx6�?t           P�@                          /�? Y�5�n?U           ��@������������������������       �        Q           p�@                         ��v�?r�q��?             @������������������������       �                     �?������������������������       �                     @                        �.w�?�<ݚ�?             K@                         �n�?���!pc�?             &@                        P-H�?z�G�z�?             $@������������������������       �                     @                        P���?�q�q�?             @                        �IN�?�q�q�?             @������������������������       �                     �?                         ��xڿ      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?       )                  ��?�ʈD��?            �E@                         ���?(N:!���?            �A@������������������������       �                     4@!       (                   f��?������?             .@"       #                  Pϕٿ8�Z$���?             *@������������������������       �                     �?$       %                 �2�?�8��8��?             (@������������������������       �                     @&       '                  s0ӿr�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @+       ,                 �̀⿨e����?            �C@������������������������       �                     &@-       4                  �$���>4և��?             <@.       3                  0mp@�eP*L��?             &@/       2                  @���?����X�?             @0       1                  ��W�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     1@6       G                  ���?��#���?�            @p@7       :                  `
ڿ0�z��?�?�             o@8       9                  �Bڿ@-�_ .�?            �B@������������������������       �                    �A@������������������������       �                      @;       F                  ��?@�� s:�?�            `j@<       =                 �Hd�? �ׁsF�?�             i@������������������������       �        x             g@>       ?                 @���?�r����?             .@������������������������       �                     �?@       E                  Έ�?@4և���?
             ,@A       D                  @ &̿r�q��?             @B       C                  SW�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �        	             &@H       K                  ��?�q�q�?
             (@I       J                 ��ſ���|���?	             &@������������������������       �                     @������������������������       �                     @������������������������       �                     �?M       �                 pʩ�?��=b4��?Q	           p�@N       �                 @���?�,���?M           Р@O       �                  �RO�?4�F��;�?           �@P       k                  ��x���B��?�           8�@Q       j                 ����*T7��?V            @_@R       _                 �/迄�����?U            �^@S       \                  `@�¿4��?�?%             J@T       U                   ��ٿ���.�6�?              G@������������������������       �        
             0@V       W                  �#�ٿףp=
�?             >@������������������������       �                     �?X       [                 P�n� 	��p�?             =@Y       Z                  �=�ؿ�����H�?             2@������������������������       ��q�q�?             @������������������������       ���S�ۿ?             .@������������������������       �                     &@]       ^                   e����q�q�?             @������������������������       �                      @������������������������       �                     @`       a                  @�ۿv���EO�?0            �Q@������������������������       �                      @b       c                 ��)��b��-8�?+            �O@������������������������       �                     @d       i                 `��翐������?)             N@e       f                  ���ڿt�F�}�?$            �I@������������������������       �                      @g       h                  ��� \� ���?#            �H@������������������������       ���[�p�?"            �G@������������������������       �                      @������������������������       �                     "@������������������������       �                      @l       �                  ��?d��n(�?�           D�@m       p                  д�ۿ�S1�<�?D           ��@n       o                 y5��q�q�?             @������������������������       �                     �?������������������������       �                      @q       r                  �:ۿP�F3���?A           ��@������������������������       �                     G@s       t                  �J7ۿ�'r�?*           (�@������������������������       �                     �?u       z                  �Eڿ��P���?)            �@v       w                 Э��|�38���?\            �d@������������������������       �                     *@x       y                 D�濪i����?V             c@������������������������       �      �?              @������������������������       �~X�<]�?R             b@{       ~                 �5�D��U��?�           ��@|       }                  qs㿠S	���?           `z@������������������������       ��/5mvq�?�             s@������������������������       �Xc!J�ƴ?H            �]@       �                 0{�߿�/FT�U�?�            �s@������������������������       �X�Cc�?             E@������������������������       �@��ɨ�?�            �p@������������������������       �        ?            �V@�       �                 `^���ϰ�T�??           `@������������������������       �        �            �o@�       �                  ��?��'�`�?�             o@������������������������       �        �            �n@������������������������       �                     @�       �                   �ۿp�,�V��?5           @~@������������������������       �                      @�       �                  ��?`��A*-�?4            ~@�       �                  p�ۿ �й���?           `{@�       �                  ��3ۿ�q�q�?             8@�       �                  0x\ۿP���Q�?             4@������������������������       �                     ,@�       �                 ���r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                  @�ڿ ��LY�s?           �y@�       �                 P�=߿h�����?             <@������������������������       �                     1@�       �                  ��ڿ�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �        �             x@������������������������       �                     F@�       �                  ��? 1�ǿ��?           @�@������������������������       �        �           ��@�       �                 P�'�?�<ݚ�?             2@�       �                  �g�ڿ      �?
             0@������������������������       �                      @������������������������       �        	             ,@������������������������       �                      @�t�b�G
      h~h,h/K ��h1��R�(KK�KK��hJ�B
       "�@     ^�@     �@     �Y@     �V@      L@     �U@              @      L@      �?      L@              L@      �?              @             0�@     �G@     h�@      B@     �@      *@     ��@      �?     p�@              @      �?              �?      @              E@      (@      @       @       @       @              @       @      @       @      �?      �?              �?      �?              �?      �?                      @      �?             �C@      @      ?@      @      4@              &@      @      &@       @              �?      &@      �?      @              @      �?      @                      �?               @       @              0@      7@      &@              @      7@      @      @      @       @      �?       @      �?                       @      @                      @              1@      o@      &@     �n@      @     �A@       @     �A@                       @      j@       @     �h@       @      g@              *@       @              �?      *@      �?      @      �?       @      �?       @                      �?      @               @              &@              @      @      @      @      @                      @      �?             ��@     ��@     ��@     0�@     �@     ��@     �@     `a@     @Y@      8@     @Y@      6@     �G@      @     �E@      @      0@              ;@      @              �?      ;@       @      0@       @       @      �?      ,@      �?      &@              @       @               @      @              K@      1@       @              G@      1@              @      G@      ,@     �B@      ,@               @     �B@      (@     �B@      $@               @      "@                       @     ��@     �\@     �@     �\@      �?       @      �?                       @     �@     @\@      G@             ��@     @\@              �?     ��@      \@      a@      =@      *@             �^@      =@      @      @     �]@      9@     `�@     �T@      x@      B@     q@      ?@     @\@      @     �p@     �G@      ;@      .@     �m@      @@     �V@              @     0@             �o@      @     �n@             �n@      @             �}@       @               @     �}@      @      {@      @      3@      @      3@      �?      ,@              @      �?              �?      @                      @     �y@      �?      ;@      �?      1@              $@      �?      $@                      �?      x@              F@              ,@     �@             ��@      ,@      @      ,@       @               @      ,@                       @�t�bubhhubehhub.