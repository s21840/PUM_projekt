��\      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �min_impurity_split�N�class_weight�N�	ccp_alpha�G        �n_features_in_�K�n_features_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�h�scalar���h'C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h'�C       �t�bK��R�}�(h	K�
node_count�KO�nodes�hhK ��h��R�(KKO��h$�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hJh'K ��hKh'K��hLh'K��hMh$�f8�����R�(Kh(NNNJ����J����K t�bK��hNhXK ��hOh'K(��hPhXK0��uK8KKt�b�BH         (                  ;ӷ?x��!���?�           ��@                         `zR�?	�h�E�?|           ��@                        ���Oi����?L	           ��@������������������������       �                   ��@                        @���?.��Ŷ�?<           �@                        �֜�?�w ��?`           ��@       
                  m�?���k4��?�           ؏@       	                 ����?���
�?�           h�@������������������������       �Ԛ܉��?�           `�@������������������������       �                     �?������������������������       �                     ,@������������������������       �        e            @Y@                         P2%ܿ�㮸DP�?�           �}@                         �jۿ�Xr��?7            �K@                         ���ܿ��:�E�?&             C@������������������������       �                      @������������������������       �
����3�?             >@������������������������       �                     1@������������������������       �        �           Pz@       #                 @���?X R&ڻ�?0           ��@                         ��ʡ)�Ŧ�?           p�@                         ��	@���"�T�?             7@                         P��?���?             4@                        �=�      �?              @������������������������       �                     �?������������������������       �                     �?                        �J��9>���?             2@������������������������       �                     ,@������������������������       ��c�����?             @                        ����|%��b�?             @������������������������       �                     �?������������������������       �                      @!       "                 �֜�?�����?�           p@������������������������       �        �           @������������������������       �                     @$       '                 �^���e���?"             A@%       &                 �I
�V�T����?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     <@)       D                 ���dԔ���?D           �@*       5                  ��'ܿZ۠�x��?�            @h@+       .                 @���?�p����?G            �Q@,       -                 �֜�?I�t���?B            �P@������������������������       �        A            @P@������������������������       �                     �?/       0                 ����?��&��?             @������������������������       �                     �?1       4                  p_�ܿ�c�����?             @2       3                   zݿ      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @6       C                  `��?����?{            �^@7       >                 P�#�?E��G9�?Y            @V@8       ;                 @���?�n$����?             >@9       :                 ���?M�)9��?             2@������������������������       �                     �?������������������������       ��S����?             1@<       =                  හ�?      �?             (@������������������������       ���&��?
             $@������������������������       �                      @?       @                  P3%ӿ�W�X�V�?;            �M@������������������������       �        !            �@@A       B                  �Hi̿���q"
�?             :@������������������������       ���&��?             @������������������������       �                     5@������������������������       �        "             A@E       F                 �֜�?4KO�?�           �@������������������������       �        h           ��@G       N                  �h.�?��M����?             :@H       M                  �3�ؿ~��kp��?             1@I       J                 ��?      �?             @������������������������       �                      @K       L                 ��+@�c�����?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �        	             "@�t�b�values�hhK ��h��R�(KKOKK��hX�B�       ��@     ΢@     �@      �@     |�@     �a@     ��@             ��@     �a@     ؎@     �`@     ��@     �`@     @�@     �`@     @�@     �`@              �?      ,@             @Y@             0}@      "@      G@      "@      =@      "@       @              5@      "@      1@             Pz@              M@     `@      9@     P@      3@      @      2@       @      �?      �?              �?      �?              1@      �?      ,@              @      �?      �?       @      �?                       @      @     @             @      @             �@@      �?      @      �?      @                      �?      <@             @X@     ��@     �T@     �[@      @     �P@      �?     @P@             @P@      �?              @       @              �?      @      �?      �?      �?      �?                      �?       @             �S@      F@     �S@      $@      6@       @      0@       @              �?      0@      �?      @      @      @      @       @             �L@       @     �@@              8@       @      @       @      5@                      A@      ,@     Й@             ��@      ,@      (@      ,@      @      @      @       @              �?      @              @      �?              &@                      "@�t�bub�_sklearn_version��0.24.2�ub.